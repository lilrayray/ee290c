module r4icLUT(
    input [10:0] io_ina,
    input [2:0] io_inb,
    output[2:0] io_r4IC
);

  wire[2:0] T0;
  wire[1:0] T1;
  reg [1:0] T2 [5119:0];
  wire[12:0] T3;
  wire[13:0] T4;
  wire[13:0] T5;
  wire[13:0] index;


  assign io_r4IC = T0;
  assign T0 = {1'h0, T1};
`ifndef SYNTHESIS
  assign T1 = T3 >= 13'h1400 ? {1{$random}} : T2[T3];
`else
  assign T1 = T2[T3];
`endif
  always @(*) begin
    T2[0] = 2'h0;
    T2[1] = 2'h0;
    T2[2] = 2'h0;
    T2[3] = 2'h0;
    T2[4] = 2'h0;
    T2[5] = 2'h1;
    T2[6] = 2'h0;
    T2[7] = 2'h0;
    T2[8] = 2'h0;
    T2[9] = 2'h0;
    T2[10] = 2'h2;
    T2[11] = 2'h0;
    T2[12] = 2'h0;
    T2[13] = 2'h0;
    T2[14] = 2'h0;
    T2[15] = 2'h3;
    T2[16] = 2'h0;
    T2[17] = 2'h0;
    T2[18] = 2'h0;
    T2[19] = 2'h0;
    T2[20] = 2'h0;
    T2[21] = 2'h1;
    T2[22] = 2'h0;
    T2[23] = 2'h0;
    T2[24] = 2'h0;
    T2[25] = 2'h1;
    T2[26] = 2'h1;
    T2[27] = 2'h0;
    T2[28] = 2'h0;
    T2[29] = 2'h0;
    T2[30] = 2'h2;
    T2[31] = 2'h1;
    T2[32] = 2'h0;
    T2[33] = 2'h0;
    T2[34] = 2'h0;
    T2[35] = 2'h3;
    T2[36] = 2'h1;
    T2[37] = 2'h0;
    T2[38] = 2'h0;
    T2[39] = 2'h0;
    T2[40] = 2'h0;
    T2[41] = 2'h2;
    T2[42] = 2'h0;
    T2[43] = 2'h0;
    T2[44] = 2'h0;
    T2[45] = 2'h1;
    T2[46] = 2'h2;
    T2[47] = 2'h0;
    T2[48] = 2'h0;
    T2[49] = 2'h0;
    T2[50] = 2'h2;
    T2[51] = 2'h2;
    T2[52] = 2'h0;
    T2[53] = 2'h0;
    T2[54] = 2'h0;
    T2[55] = 2'h3;
    T2[56] = 2'h2;
    T2[57] = 2'h0;
    T2[58] = 2'h0;
    T2[59] = 2'h0;
    T2[60] = 2'h0;
    T2[61] = 2'h3;
    T2[62] = 2'h0;
    T2[63] = 2'h0;
    T2[64] = 2'h0;
    T2[65] = 2'h1;
    T2[66] = 2'h3;
    T2[67] = 2'h0;
    T2[68] = 2'h0;
    T2[69] = 2'h0;
    T2[70] = 2'h2;
    T2[71] = 2'h3;
    T2[72] = 2'h0;
    T2[73] = 2'h0;
    T2[74] = 2'h0;
    T2[75] = 2'h3;
    T2[76] = 2'h3;
    T2[77] = 2'h0;
    T2[78] = 2'h0;
    T2[79] = 2'h0;
    T2[80] = 2'h0;
    T2[81] = 2'h0;
    T2[82] = 2'h1;
    T2[83] = 2'h0;
    T2[84] = 2'h0;
    T2[85] = 2'h1;
    T2[86] = 2'h0;
    T2[87] = 2'h1;
    T2[88] = 2'h0;
    T2[89] = 2'h0;
    T2[90] = 2'h2;
    T2[91] = 2'h0;
    T2[92] = 2'h1;
    T2[93] = 2'h0;
    T2[94] = 2'h0;
    T2[95] = 2'h3;
    T2[96] = 2'h0;
    T2[97] = 2'h1;
    T2[98] = 2'h0;
    T2[99] = 2'h0;
    T2[100] = 2'h0;
    T2[101] = 2'h1;
    T2[102] = 2'h1;
    T2[103] = 2'h0;
    T2[104] = 2'h0;
    T2[105] = 2'h1;
    T2[106] = 2'h1;
    T2[107] = 2'h1;
    T2[108] = 2'h0;
    T2[109] = 2'h0;
    T2[110] = 2'h2;
    T2[111] = 2'h1;
    T2[112] = 2'h1;
    T2[113] = 2'h0;
    T2[114] = 2'h0;
    T2[115] = 2'h3;
    T2[116] = 2'h1;
    T2[117] = 2'h1;
    T2[118] = 2'h0;
    T2[119] = 2'h0;
    T2[120] = 2'h0;
    T2[121] = 2'h2;
    T2[122] = 2'h1;
    T2[123] = 2'h0;
    T2[124] = 2'h0;
    T2[125] = 2'h1;
    T2[126] = 2'h2;
    T2[127] = 2'h1;
    T2[128] = 2'h0;
    T2[129] = 2'h0;
    T2[130] = 2'h2;
    T2[131] = 2'h2;
    T2[132] = 2'h1;
    T2[133] = 2'h0;
    T2[134] = 2'h0;
    T2[135] = 2'h3;
    T2[136] = 2'h2;
    T2[137] = 2'h1;
    T2[138] = 2'h0;
    T2[139] = 2'h0;
    T2[140] = 2'h0;
    T2[141] = 2'h3;
    T2[142] = 2'h1;
    T2[143] = 2'h0;
    T2[144] = 2'h0;
    T2[145] = 2'h1;
    T2[146] = 2'h3;
    T2[147] = 2'h1;
    T2[148] = 2'h0;
    T2[149] = 2'h0;
    T2[150] = 2'h2;
    T2[151] = 2'h3;
    T2[152] = 2'h1;
    T2[153] = 2'h0;
    T2[154] = 2'h0;
    T2[155] = 2'h3;
    T2[156] = 2'h3;
    T2[157] = 2'h1;
    T2[158] = 2'h0;
    T2[159] = 2'h0;
    T2[160] = 2'h0;
    T2[161] = 2'h0;
    T2[162] = 2'h2;
    T2[163] = 2'h0;
    T2[164] = 2'h0;
    T2[165] = 2'h1;
    T2[166] = 2'h0;
    T2[167] = 2'h2;
    T2[168] = 2'h0;
    T2[169] = 2'h0;
    T2[170] = 2'h2;
    T2[171] = 2'h0;
    T2[172] = 2'h2;
    T2[173] = 2'h0;
    T2[174] = 2'h0;
    T2[175] = 2'h3;
    T2[176] = 2'h0;
    T2[177] = 2'h2;
    T2[178] = 2'h0;
    T2[179] = 2'h0;
    T2[180] = 2'h0;
    T2[181] = 2'h1;
    T2[182] = 2'h2;
    T2[183] = 2'h0;
    T2[184] = 2'h0;
    T2[185] = 2'h1;
    T2[186] = 2'h1;
    T2[187] = 2'h2;
    T2[188] = 2'h0;
    T2[189] = 2'h0;
    T2[190] = 2'h2;
    T2[191] = 2'h1;
    T2[192] = 2'h2;
    T2[193] = 2'h0;
    T2[194] = 2'h0;
    T2[195] = 2'h3;
    T2[196] = 2'h1;
    T2[197] = 2'h2;
    T2[198] = 2'h0;
    T2[199] = 2'h0;
    T2[200] = 2'h0;
    T2[201] = 2'h2;
    T2[202] = 2'h2;
    T2[203] = 2'h0;
    T2[204] = 2'h0;
    T2[205] = 2'h1;
    T2[206] = 2'h2;
    T2[207] = 2'h2;
    T2[208] = 2'h0;
    T2[209] = 2'h0;
    T2[210] = 2'h2;
    T2[211] = 2'h2;
    T2[212] = 2'h2;
    T2[213] = 2'h0;
    T2[214] = 2'h0;
    T2[215] = 2'h3;
    T2[216] = 2'h2;
    T2[217] = 2'h2;
    T2[218] = 2'h0;
    T2[219] = 2'h0;
    T2[220] = 2'h0;
    T2[221] = 2'h3;
    T2[222] = 2'h2;
    T2[223] = 2'h0;
    T2[224] = 2'h0;
    T2[225] = 2'h1;
    T2[226] = 2'h3;
    T2[227] = 2'h2;
    T2[228] = 2'h0;
    T2[229] = 2'h0;
    T2[230] = 2'h2;
    T2[231] = 2'h3;
    T2[232] = 2'h2;
    T2[233] = 2'h0;
    T2[234] = 2'h0;
    T2[235] = 2'h3;
    T2[236] = 2'h3;
    T2[237] = 2'h2;
    T2[238] = 2'h0;
    T2[239] = 2'h0;
    T2[240] = 2'h0;
    T2[241] = 2'h0;
    T2[242] = 2'h3;
    T2[243] = 2'h0;
    T2[244] = 2'h0;
    T2[245] = 2'h1;
    T2[246] = 2'h0;
    T2[247] = 2'h3;
    T2[248] = 2'h0;
    T2[249] = 2'h0;
    T2[250] = 2'h2;
    T2[251] = 2'h0;
    T2[252] = 2'h3;
    T2[253] = 2'h0;
    T2[254] = 2'h0;
    T2[255] = 2'h3;
    T2[256] = 2'h0;
    T2[257] = 2'h3;
    T2[258] = 2'h0;
    T2[259] = 2'h0;
    T2[260] = 2'h0;
    T2[261] = 2'h1;
    T2[262] = 2'h3;
    T2[263] = 2'h0;
    T2[264] = 2'h0;
    T2[265] = 2'h1;
    T2[266] = 2'h1;
    T2[267] = 2'h3;
    T2[268] = 2'h0;
    T2[269] = 2'h0;
    T2[270] = 2'h2;
    T2[271] = 2'h1;
    T2[272] = 2'h3;
    T2[273] = 2'h0;
    T2[274] = 2'h0;
    T2[275] = 2'h3;
    T2[276] = 2'h1;
    T2[277] = 2'h3;
    T2[278] = 2'h0;
    T2[279] = 2'h0;
    T2[280] = 2'h0;
    T2[281] = 2'h2;
    T2[282] = 2'h3;
    T2[283] = 2'h0;
    T2[284] = 2'h0;
    T2[285] = 2'h1;
    T2[286] = 2'h2;
    T2[287] = 2'h3;
    T2[288] = 2'h0;
    T2[289] = 2'h0;
    T2[290] = 2'h2;
    T2[291] = 2'h2;
    T2[292] = 2'h3;
    T2[293] = 2'h0;
    T2[294] = 2'h0;
    T2[295] = 2'h3;
    T2[296] = 2'h2;
    T2[297] = 2'h3;
    T2[298] = 2'h0;
    T2[299] = 2'h0;
    T2[300] = 2'h0;
    T2[301] = 2'h3;
    T2[302] = 2'h3;
    T2[303] = 2'h0;
    T2[304] = 2'h0;
    T2[305] = 2'h1;
    T2[306] = 2'h3;
    T2[307] = 2'h3;
    T2[308] = 2'h0;
    T2[309] = 2'h0;
    T2[310] = 2'h2;
    T2[311] = 2'h3;
    T2[312] = 2'h3;
    T2[313] = 2'h0;
    T2[314] = 2'h0;
    T2[315] = 2'h3;
    T2[316] = 2'h3;
    T2[317] = 2'h3;
    T2[318] = 2'h0;
    T2[319] = 2'h0;
    T2[320] = 2'h0;
    T2[321] = 2'h0;
    T2[322] = 2'h0;
    T2[323] = 2'h1;
    T2[324] = 2'h0;
    T2[325] = 2'h1;
    T2[326] = 2'h0;
    T2[327] = 2'h0;
    T2[328] = 2'h1;
    T2[329] = 2'h0;
    T2[330] = 2'h2;
    T2[331] = 2'h0;
    T2[332] = 2'h0;
    T2[333] = 2'h1;
    T2[334] = 2'h0;
    T2[335] = 2'h3;
    T2[336] = 2'h0;
    T2[337] = 2'h0;
    T2[338] = 2'h1;
    T2[339] = 2'h0;
    T2[340] = 2'h0;
    T2[341] = 2'h1;
    T2[342] = 2'h0;
    T2[343] = 2'h1;
    T2[344] = 2'h0;
    T2[345] = 2'h1;
    T2[346] = 2'h1;
    T2[347] = 2'h0;
    T2[348] = 2'h1;
    T2[349] = 2'h0;
    T2[350] = 2'h2;
    T2[351] = 2'h1;
    T2[352] = 2'h0;
    T2[353] = 2'h1;
    T2[354] = 2'h0;
    T2[355] = 2'h3;
    T2[356] = 2'h1;
    T2[357] = 2'h0;
    T2[358] = 2'h1;
    T2[359] = 2'h0;
    T2[360] = 2'h0;
    T2[361] = 2'h2;
    T2[362] = 2'h0;
    T2[363] = 2'h1;
    T2[364] = 2'h0;
    T2[365] = 2'h1;
    T2[366] = 2'h2;
    T2[367] = 2'h0;
    T2[368] = 2'h1;
    T2[369] = 2'h0;
    T2[370] = 2'h2;
    T2[371] = 2'h2;
    T2[372] = 2'h0;
    T2[373] = 2'h1;
    T2[374] = 2'h0;
    T2[375] = 2'h3;
    T2[376] = 2'h2;
    T2[377] = 2'h0;
    T2[378] = 2'h1;
    T2[379] = 2'h0;
    T2[380] = 2'h0;
    T2[381] = 2'h3;
    T2[382] = 2'h0;
    T2[383] = 2'h1;
    T2[384] = 2'h0;
    T2[385] = 2'h1;
    T2[386] = 2'h3;
    T2[387] = 2'h0;
    T2[388] = 2'h1;
    T2[389] = 2'h0;
    T2[390] = 2'h2;
    T2[391] = 2'h3;
    T2[392] = 2'h0;
    T2[393] = 2'h1;
    T2[394] = 2'h0;
    T2[395] = 2'h3;
    T2[396] = 2'h3;
    T2[397] = 2'h0;
    T2[398] = 2'h1;
    T2[399] = 2'h0;
    T2[400] = 2'h0;
    T2[401] = 2'h0;
    T2[402] = 2'h1;
    T2[403] = 2'h1;
    T2[404] = 2'h0;
    T2[405] = 2'h1;
    T2[406] = 2'h0;
    T2[407] = 2'h1;
    T2[408] = 2'h1;
    T2[409] = 2'h0;
    T2[410] = 2'h2;
    T2[411] = 2'h0;
    T2[412] = 2'h1;
    T2[413] = 2'h1;
    T2[414] = 2'h0;
    T2[415] = 2'h3;
    T2[416] = 2'h0;
    T2[417] = 2'h1;
    T2[418] = 2'h1;
    T2[419] = 2'h0;
    T2[420] = 2'h0;
    T2[421] = 2'h1;
    T2[422] = 2'h1;
    T2[423] = 2'h1;
    T2[424] = 2'h0;
    T2[425] = 2'h1;
    T2[426] = 2'h1;
    T2[427] = 2'h1;
    T2[428] = 2'h1;
    T2[429] = 2'h0;
    T2[430] = 2'h2;
    T2[431] = 2'h1;
    T2[432] = 2'h1;
    T2[433] = 2'h1;
    T2[434] = 2'h0;
    T2[435] = 2'h3;
    T2[436] = 2'h1;
    T2[437] = 2'h1;
    T2[438] = 2'h1;
    T2[439] = 2'h0;
    T2[440] = 2'h0;
    T2[441] = 2'h2;
    T2[442] = 2'h1;
    T2[443] = 2'h1;
    T2[444] = 2'h0;
    T2[445] = 2'h1;
    T2[446] = 2'h2;
    T2[447] = 2'h1;
    T2[448] = 2'h1;
    T2[449] = 2'h0;
    T2[450] = 2'h2;
    T2[451] = 2'h2;
    T2[452] = 2'h1;
    T2[453] = 2'h1;
    T2[454] = 2'h0;
    T2[455] = 2'h3;
    T2[456] = 2'h2;
    T2[457] = 2'h1;
    T2[458] = 2'h1;
    T2[459] = 2'h0;
    T2[460] = 2'h0;
    T2[461] = 2'h3;
    T2[462] = 2'h1;
    T2[463] = 2'h1;
    T2[464] = 2'h0;
    T2[465] = 2'h1;
    T2[466] = 2'h3;
    T2[467] = 2'h1;
    T2[468] = 2'h1;
    T2[469] = 2'h0;
    T2[470] = 2'h2;
    T2[471] = 2'h3;
    T2[472] = 2'h1;
    T2[473] = 2'h1;
    T2[474] = 2'h0;
    T2[475] = 2'h3;
    T2[476] = 2'h3;
    T2[477] = 2'h1;
    T2[478] = 2'h1;
    T2[479] = 2'h0;
    T2[480] = 2'h0;
    T2[481] = 2'h0;
    T2[482] = 2'h2;
    T2[483] = 2'h1;
    T2[484] = 2'h0;
    T2[485] = 2'h1;
    T2[486] = 2'h0;
    T2[487] = 2'h2;
    T2[488] = 2'h1;
    T2[489] = 2'h0;
    T2[490] = 2'h2;
    T2[491] = 2'h0;
    T2[492] = 2'h2;
    T2[493] = 2'h1;
    T2[494] = 2'h0;
    T2[495] = 2'h3;
    T2[496] = 2'h0;
    T2[497] = 2'h2;
    T2[498] = 2'h1;
    T2[499] = 2'h0;
    T2[500] = 2'h0;
    T2[501] = 2'h1;
    T2[502] = 2'h2;
    T2[503] = 2'h1;
    T2[504] = 2'h0;
    T2[505] = 2'h1;
    T2[506] = 2'h1;
    T2[507] = 2'h2;
    T2[508] = 2'h1;
    T2[509] = 2'h0;
    T2[510] = 2'h2;
    T2[511] = 2'h1;
    T2[512] = 2'h2;
    T2[513] = 2'h1;
    T2[514] = 2'h0;
    T2[515] = 2'h3;
    T2[516] = 2'h1;
    T2[517] = 2'h2;
    T2[518] = 2'h1;
    T2[519] = 2'h0;
    T2[520] = 2'h0;
    T2[521] = 2'h2;
    T2[522] = 2'h2;
    T2[523] = 2'h1;
    T2[524] = 2'h0;
    T2[525] = 2'h1;
    T2[526] = 2'h2;
    T2[527] = 2'h2;
    T2[528] = 2'h1;
    T2[529] = 2'h0;
    T2[530] = 2'h2;
    T2[531] = 2'h2;
    T2[532] = 2'h2;
    T2[533] = 2'h1;
    T2[534] = 2'h0;
    T2[535] = 2'h3;
    T2[536] = 2'h2;
    T2[537] = 2'h2;
    T2[538] = 2'h1;
    T2[539] = 2'h0;
    T2[540] = 2'h0;
    T2[541] = 2'h3;
    T2[542] = 2'h2;
    T2[543] = 2'h1;
    T2[544] = 2'h0;
    T2[545] = 2'h1;
    T2[546] = 2'h3;
    T2[547] = 2'h2;
    T2[548] = 2'h1;
    T2[549] = 2'h0;
    T2[550] = 2'h2;
    T2[551] = 2'h3;
    T2[552] = 2'h2;
    T2[553] = 2'h1;
    T2[554] = 2'h0;
    T2[555] = 2'h3;
    T2[556] = 2'h3;
    T2[557] = 2'h2;
    T2[558] = 2'h1;
    T2[559] = 2'h0;
    T2[560] = 2'h0;
    T2[561] = 2'h0;
    T2[562] = 2'h3;
    T2[563] = 2'h1;
    T2[564] = 2'h0;
    T2[565] = 2'h1;
    T2[566] = 2'h0;
    T2[567] = 2'h3;
    T2[568] = 2'h1;
    T2[569] = 2'h0;
    T2[570] = 2'h2;
    T2[571] = 2'h0;
    T2[572] = 2'h3;
    T2[573] = 2'h1;
    T2[574] = 2'h0;
    T2[575] = 2'h3;
    T2[576] = 2'h0;
    T2[577] = 2'h3;
    T2[578] = 2'h1;
    T2[579] = 2'h0;
    T2[580] = 2'h0;
    T2[581] = 2'h1;
    T2[582] = 2'h3;
    T2[583] = 2'h1;
    T2[584] = 2'h0;
    T2[585] = 2'h1;
    T2[586] = 2'h1;
    T2[587] = 2'h3;
    T2[588] = 2'h1;
    T2[589] = 2'h0;
    T2[590] = 2'h2;
    T2[591] = 2'h1;
    T2[592] = 2'h3;
    T2[593] = 2'h1;
    T2[594] = 2'h0;
    T2[595] = 2'h3;
    T2[596] = 2'h1;
    T2[597] = 2'h3;
    T2[598] = 2'h1;
    T2[599] = 2'h0;
    T2[600] = 2'h0;
    T2[601] = 2'h2;
    T2[602] = 2'h3;
    T2[603] = 2'h1;
    T2[604] = 2'h0;
    T2[605] = 2'h1;
    T2[606] = 2'h2;
    T2[607] = 2'h3;
    T2[608] = 2'h1;
    T2[609] = 2'h0;
    T2[610] = 2'h2;
    T2[611] = 2'h2;
    T2[612] = 2'h3;
    T2[613] = 2'h1;
    T2[614] = 2'h0;
    T2[615] = 2'h3;
    T2[616] = 2'h2;
    T2[617] = 2'h3;
    T2[618] = 2'h1;
    T2[619] = 2'h0;
    T2[620] = 2'h0;
    T2[621] = 2'h3;
    T2[622] = 2'h3;
    T2[623] = 2'h1;
    T2[624] = 2'h0;
    T2[625] = 2'h1;
    T2[626] = 2'h3;
    T2[627] = 2'h3;
    T2[628] = 2'h1;
    T2[629] = 2'h0;
    T2[630] = 2'h2;
    T2[631] = 2'h3;
    T2[632] = 2'h3;
    T2[633] = 2'h1;
    T2[634] = 2'h0;
    T2[635] = 2'h3;
    T2[636] = 2'h3;
    T2[637] = 2'h3;
    T2[638] = 2'h1;
    T2[639] = 2'h0;
    T2[640] = 2'h0;
    T2[641] = 2'h0;
    T2[642] = 2'h0;
    T2[643] = 2'h2;
    T2[644] = 2'h0;
    T2[645] = 2'h1;
    T2[646] = 2'h0;
    T2[647] = 2'h0;
    T2[648] = 2'h2;
    T2[649] = 2'h0;
    T2[650] = 2'h2;
    T2[651] = 2'h0;
    T2[652] = 2'h0;
    T2[653] = 2'h2;
    T2[654] = 2'h0;
    T2[655] = 2'h3;
    T2[656] = 2'h0;
    T2[657] = 2'h0;
    T2[658] = 2'h2;
    T2[659] = 2'h0;
    T2[660] = 2'h0;
    T2[661] = 2'h1;
    T2[662] = 2'h0;
    T2[663] = 2'h2;
    T2[664] = 2'h0;
    T2[665] = 2'h1;
    T2[666] = 2'h1;
    T2[667] = 2'h0;
    T2[668] = 2'h2;
    T2[669] = 2'h0;
    T2[670] = 2'h2;
    T2[671] = 2'h1;
    T2[672] = 2'h0;
    T2[673] = 2'h2;
    T2[674] = 2'h0;
    T2[675] = 2'h3;
    T2[676] = 2'h1;
    T2[677] = 2'h0;
    T2[678] = 2'h2;
    T2[679] = 2'h0;
    T2[680] = 2'h0;
    T2[681] = 2'h2;
    T2[682] = 2'h0;
    T2[683] = 2'h2;
    T2[684] = 2'h0;
    T2[685] = 2'h1;
    T2[686] = 2'h2;
    T2[687] = 2'h0;
    T2[688] = 2'h2;
    T2[689] = 2'h0;
    T2[690] = 2'h2;
    T2[691] = 2'h2;
    T2[692] = 2'h0;
    T2[693] = 2'h2;
    T2[694] = 2'h0;
    T2[695] = 2'h3;
    T2[696] = 2'h2;
    T2[697] = 2'h0;
    T2[698] = 2'h2;
    T2[699] = 2'h0;
    T2[700] = 2'h0;
    T2[701] = 2'h3;
    T2[702] = 2'h0;
    T2[703] = 2'h2;
    T2[704] = 2'h0;
    T2[705] = 2'h1;
    T2[706] = 2'h3;
    T2[707] = 2'h0;
    T2[708] = 2'h2;
    T2[709] = 2'h0;
    T2[710] = 2'h2;
    T2[711] = 2'h3;
    T2[712] = 2'h0;
    T2[713] = 2'h2;
    T2[714] = 2'h0;
    T2[715] = 2'h3;
    T2[716] = 2'h3;
    T2[717] = 2'h0;
    T2[718] = 2'h2;
    T2[719] = 2'h0;
    T2[720] = 2'h0;
    T2[721] = 2'h0;
    T2[722] = 2'h1;
    T2[723] = 2'h2;
    T2[724] = 2'h0;
    T2[725] = 2'h1;
    T2[726] = 2'h0;
    T2[727] = 2'h1;
    T2[728] = 2'h2;
    T2[729] = 2'h0;
    T2[730] = 2'h2;
    T2[731] = 2'h0;
    T2[732] = 2'h1;
    T2[733] = 2'h2;
    T2[734] = 2'h0;
    T2[735] = 2'h3;
    T2[736] = 2'h0;
    T2[737] = 2'h1;
    T2[738] = 2'h2;
    T2[739] = 2'h0;
    T2[740] = 2'h0;
    T2[741] = 2'h1;
    T2[742] = 2'h1;
    T2[743] = 2'h2;
    T2[744] = 2'h0;
    T2[745] = 2'h1;
    T2[746] = 2'h1;
    T2[747] = 2'h1;
    T2[748] = 2'h2;
    T2[749] = 2'h0;
    T2[750] = 2'h2;
    T2[751] = 2'h1;
    T2[752] = 2'h1;
    T2[753] = 2'h2;
    T2[754] = 2'h0;
    T2[755] = 2'h3;
    T2[756] = 2'h1;
    T2[757] = 2'h1;
    T2[758] = 2'h2;
    T2[759] = 2'h0;
    T2[760] = 2'h0;
    T2[761] = 2'h2;
    T2[762] = 2'h1;
    T2[763] = 2'h2;
    T2[764] = 2'h0;
    T2[765] = 2'h1;
    T2[766] = 2'h2;
    T2[767] = 2'h1;
    T2[768] = 2'h2;
    T2[769] = 2'h0;
    T2[770] = 2'h2;
    T2[771] = 2'h2;
    T2[772] = 2'h1;
    T2[773] = 2'h2;
    T2[774] = 2'h0;
    T2[775] = 2'h3;
    T2[776] = 2'h2;
    T2[777] = 2'h1;
    T2[778] = 2'h2;
    T2[779] = 2'h0;
    T2[780] = 2'h0;
    T2[781] = 2'h3;
    T2[782] = 2'h1;
    T2[783] = 2'h2;
    T2[784] = 2'h0;
    T2[785] = 2'h1;
    T2[786] = 2'h3;
    T2[787] = 2'h1;
    T2[788] = 2'h2;
    T2[789] = 2'h0;
    T2[790] = 2'h2;
    T2[791] = 2'h3;
    T2[792] = 2'h1;
    T2[793] = 2'h2;
    T2[794] = 2'h0;
    T2[795] = 2'h3;
    T2[796] = 2'h3;
    T2[797] = 2'h1;
    T2[798] = 2'h2;
    T2[799] = 2'h0;
    T2[800] = 2'h0;
    T2[801] = 2'h0;
    T2[802] = 2'h2;
    T2[803] = 2'h2;
    T2[804] = 2'h0;
    T2[805] = 2'h1;
    T2[806] = 2'h0;
    T2[807] = 2'h2;
    T2[808] = 2'h2;
    T2[809] = 2'h0;
    T2[810] = 2'h2;
    T2[811] = 2'h0;
    T2[812] = 2'h2;
    T2[813] = 2'h2;
    T2[814] = 2'h0;
    T2[815] = 2'h3;
    T2[816] = 2'h0;
    T2[817] = 2'h2;
    T2[818] = 2'h2;
    T2[819] = 2'h0;
    T2[820] = 2'h0;
    T2[821] = 2'h1;
    T2[822] = 2'h2;
    T2[823] = 2'h2;
    T2[824] = 2'h0;
    T2[825] = 2'h1;
    T2[826] = 2'h1;
    T2[827] = 2'h2;
    T2[828] = 2'h2;
    T2[829] = 2'h0;
    T2[830] = 2'h2;
    T2[831] = 2'h1;
    T2[832] = 2'h2;
    T2[833] = 2'h2;
    T2[834] = 2'h0;
    T2[835] = 2'h3;
    T2[836] = 2'h1;
    T2[837] = 2'h2;
    T2[838] = 2'h2;
    T2[839] = 2'h0;
    T2[840] = 2'h0;
    T2[841] = 2'h2;
    T2[842] = 2'h2;
    T2[843] = 2'h2;
    T2[844] = 2'h0;
    T2[845] = 2'h1;
    T2[846] = 2'h2;
    T2[847] = 2'h2;
    T2[848] = 2'h2;
    T2[849] = 2'h0;
    T2[850] = 2'h2;
    T2[851] = 2'h2;
    T2[852] = 2'h2;
    T2[853] = 2'h2;
    T2[854] = 2'h0;
    T2[855] = 2'h3;
    T2[856] = 2'h2;
    T2[857] = 2'h2;
    T2[858] = 2'h2;
    T2[859] = 2'h0;
    T2[860] = 2'h0;
    T2[861] = 2'h3;
    T2[862] = 2'h2;
    T2[863] = 2'h2;
    T2[864] = 2'h0;
    T2[865] = 2'h1;
    T2[866] = 2'h3;
    T2[867] = 2'h2;
    T2[868] = 2'h2;
    T2[869] = 2'h0;
    T2[870] = 2'h2;
    T2[871] = 2'h3;
    T2[872] = 2'h2;
    T2[873] = 2'h2;
    T2[874] = 2'h0;
    T2[875] = 2'h3;
    T2[876] = 2'h3;
    T2[877] = 2'h2;
    T2[878] = 2'h2;
    T2[879] = 2'h0;
    T2[880] = 2'h0;
    T2[881] = 2'h0;
    T2[882] = 2'h3;
    T2[883] = 2'h2;
    T2[884] = 2'h0;
    T2[885] = 2'h1;
    T2[886] = 2'h0;
    T2[887] = 2'h3;
    T2[888] = 2'h2;
    T2[889] = 2'h0;
    T2[890] = 2'h2;
    T2[891] = 2'h0;
    T2[892] = 2'h3;
    T2[893] = 2'h2;
    T2[894] = 2'h0;
    T2[895] = 2'h3;
    T2[896] = 2'h0;
    T2[897] = 2'h3;
    T2[898] = 2'h2;
    T2[899] = 2'h0;
    T2[900] = 2'h0;
    T2[901] = 2'h1;
    T2[902] = 2'h3;
    T2[903] = 2'h2;
    T2[904] = 2'h0;
    T2[905] = 2'h1;
    T2[906] = 2'h1;
    T2[907] = 2'h3;
    T2[908] = 2'h2;
    T2[909] = 2'h0;
    T2[910] = 2'h2;
    T2[911] = 2'h1;
    T2[912] = 2'h3;
    T2[913] = 2'h2;
    T2[914] = 2'h0;
    T2[915] = 2'h3;
    T2[916] = 2'h1;
    T2[917] = 2'h3;
    T2[918] = 2'h2;
    T2[919] = 2'h0;
    T2[920] = 2'h0;
    T2[921] = 2'h2;
    T2[922] = 2'h3;
    T2[923] = 2'h2;
    T2[924] = 2'h0;
    T2[925] = 2'h1;
    T2[926] = 2'h2;
    T2[927] = 2'h3;
    T2[928] = 2'h2;
    T2[929] = 2'h0;
    T2[930] = 2'h2;
    T2[931] = 2'h2;
    T2[932] = 2'h3;
    T2[933] = 2'h2;
    T2[934] = 2'h0;
    T2[935] = 2'h3;
    T2[936] = 2'h2;
    T2[937] = 2'h3;
    T2[938] = 2'h2;
    T2[939] = 2'h0;
    T2[940] = 2'h0;
    T2[941] = 2'h3;
    T2[942] = 2'h3;
    T2[943] = 2'h2;
    T2[944] = 2'h0;
    T2[945] = 2'h1;
    T2[946] = 2'h3;
    T2[947] = 2'h3;
    T2[948] = 2'h2;
    T2[949] = 2'h0;
    T2[950] = 2'h2;
    T2[951] = 2'h3;
    T2[952] = 2'h3;
    T2[953] = 2'h2;
    T2[954] = 2'h0;
    T2[955] = 2'h3;
    T2[956] = 2'h3;
    T2[957] = 2'h3;
    T2[958] = 2'h2;
    T2[959] = 2'h0;
    T2[960] = 2'h0;
    T2[961] = 2'h0;
    T2[962] = 2'h0;
    T2[963] = 2'h3;
    T2[964] = 2'h0;
    T2[965] = 2'h1;
    T2[966] = 2'h0;
    T2[967] = 2'h0;
    T2[968] = 2'h3;
    T2[969] = 2'h0;
    T2[970] = 2'h2;
    T2[971] = 2'h0;
    T2[972] = 2'h0;
    T2[973] = 2'h3;
    T2[974] = 2'h0;
    T2[975] = 2'h3;
    T2[976] = 2'h0;
    T2[977] = 2'h0;
    T2[978] = 2'h3;
    T2[979] = 2'h0;
    T2[980] = 2'h0;
    T2[981] = 2'h1;
    T2[982] = 2'h0;
    T2[983] = 2'h3;
    T2[984] = 2'h0;
    T2[985] = 2'h1;
    T2[986] = 2'h1;
    T2[987] = 2'h0;
    T2[988] = 2'h3;
    T2[989] = 2'h0;
    T2[990] = 2'h2;
    T2[991] = 2'h1;
    T2[992] = 2'h0;
    T2[993] = 2'h3;
    T2[994] = 2'h0;
    T2[995] = 2'h3;
    T2[996] = 2'h1;
    T2[997] = 2'h0;
    T2[998] = 2'h3;
    T2[999] = 2'h0;
    T2[1000] = 2'h0;
    T2[1001] = 2'h2;
    T2[1002] = 2'h0;
    T2[1003] = 2'h3;
    T2[1004] = 2'h0;
    T2[1005] = 2'h1;
    T2[1006] = 2'h2;
    T2[1007] = 2'h0;
    T2[1008] = 2'h3;
    T2[1009] = 2'h0;
    T2[1010] = 2'h2;
    T2[1011] = 2'h2;
    T2[1012] = 2'h0;
    T2[1013] = 2'h3;
    T2[1014] = 2'h0;
    T2[1015] = 2'h3;
    T2[1016] = 2'h2;
    T2[1017] = 2'h0;
    T2[1018] = 2'h3;
    T2[1019] = 2'h0;
    T2[1020] = 2'h0;
    T2[1021] = 2'h3;
    T2[1022] = 2'h0;
    T2[1023] = 2'h3;
    T2[1024] = 2'h0;
    T2[1025] = 2'h1;
    T2[1026] = 2'h3;
    T2[1027] = 2'h0;
    T2[1028] = 2'h3;
    T2[1029] = 2'h0;
    T2[1030] = 2'h2;
    T2[1031] = 2'h3;
    T2[1032] = 2'h0;
    T2[1033] = 2'h3;
    T2[1034] = 2'h0;
    T2[1035] = 2'h3;
    T2[1036] = 2'h3;
    T2[1037] = 2'h0;
    T2[1038] = 2'h3;
    T2[1039] = 2'h0;
    T2[1040] = 2'h0;
    T2[1041] = 2'h0;
    T2[1042] = 2'h1;
    T2[1043] = 2'h3;
    T2[1044] = 2'h0;
    T2[1045] = 2'h1;
    T2[1046] = 2'h0;
    T2[1047] = 2'h1;
    T2[1048] = 2'h3;
    T2[1049] = 2'h0;
    T2[1050] = 2'h2;
    T2[1051] = 2'h0;
    T2[1052] = 2'h1;
    T2[1053] = 2'h3;
    T2[1054] = 2'h0;
    T2[1055] = 2'h3;
    T2[1056] = 2'h0;
    T2[1057] = 2'h1;
    T2[1058] = 2'h3;
    T2[1059] = 2'h0;
    T2[1060] = 2'h0;
    T2[1061] = 2'h1;
    T2[1062] = 2'h1;
    T2[1063] = 2'h3;
    T2[1064] = 2'h0;
    T2[1065] = 2'h1;
    T2[1066] = 2'h1;
    T2[1067] = 2'h1;
    T2[1068] = 2'h3;
    T2[1069] = 2'h0;
    T2[1070] = 2'h2;
    T2[1071] = 2'h1;
    T2[1072] = 2'h1;
    T2[1073] = 2'h3;
    T2[1074] = 2'h0;
    T2[1075] = 2'h3;
    T2[1076] = 2'h1;
    T2[1077] = 2'h1;
    T2[1078] = 2'h3;
    T2[1079] = 2'h0;
    T2[1080] = 2'h0;
    T2[1081] = 2'h2;
    T2[1082] = 2'h1;
    T2[1083] = 2'h3;
    T2[1084] = 2'h0;
    T2[1085] = 2'h1;
    T2[1086] = 2'h2;
    T2[1087] = 2'h1;
    T2[1088] = 2'h3;
    T2[1089] = 2'h0;
    T2[1090] = 2'h2;
    T2[1091] = 2'h2;
    T2[1092] = 2'h1;
    T2[1093] = 2'h3;
    T2[1094] = 2'h0;
    T2[1095] = 2'h3;
    T2[1096] = 2'h2;
    T2[1097] = 2'h1;
    T2[1098] = 2'h3;
    T2[1099] = 2'h0;
    T2[1100] = 2'h0;
    T2[1101] = 2'h3;
    T2[1102] = 2'h1;
    T2[1103] = 2'h3;
    T2[1104] = 2'h0;
    T2[1105] = 2'h1;
    T2[1106] = 2'h3;
    T2[1107] = 2'h1;
    T2[1108] = 2'h3;
    T2[1109] = 2'h0;
    T2[1110] = 2'h2;
    T2[1111] = 2'h3;
    T2[1112] = 2'h1;
    T2[1113] = 2'h3;
    T2[1114] = 2'h0;
    T2[1115] = 2'h3;
    T2[1116] = 2'h3;
    T2[1117] = 2'h1;
    T2[1118] = 2'h3;
    T2[1119] = 2'h0;
    T2[1120] = 2'h0;
    T2[1121] = 2'h0;
    T2[1122] = 2'h2;
    T2[1123] = 2'h3;
    T2[1124] = 2'h0;
    T2[1125] = 2'h1;
    T2[1126] = 2'h0;
    T2[1127] = 2'h2;
    T2[1128] = 2'h3;
    T2[1129] = 2'h0;
    T2[1130] = 2'h2;
    T2[1131] = 2'h0;
    T2[1132] = 2'h2;
    T2[1133] = 2'h3;
    T2[1134] = 2'h0;
    T2[1135] = 2'h3;
    T2[1136] = 2'h0;
    T2[1137] = 2'h2;
    T2[1138] = 2'h3;
    T2[1139] = 2'h0;
    T2[1140] = 2'h0;
    T2[1141] = 2'h1;
    T2[1142] = 2'h2;
    T2[1143] = 2'h3;
    T2[1144] = 2'h0;
    T2[1145] = 2'h1;
    T2[1146] = 2'h1;
    T2[1147] = 2'h2;
    T2[1148] = 2'h3;
    T2[1149] = 2'h0;
    T2[1150] = 2'h2;
    T2[1151] = 2'h1;
    T2[1152] = 2'h2;
    T2[1153] = 2'h3;
    T2[1154] = 2'h0;
    T2[1155] = 2'h3;
    T2[1156] = 2'h1;
    T2[1157] = 2'h2;
    T2[1158] = 2'h3;
    T2[1159] = 2'h0;
    T2[1160] = 2'h0;
    T2[1161] = 2'h2;
    T2[1162] = 2'h2;
    T2[1163] = 2'h3;
    T2[1164] = 2'h0;
    T2[1165] = 2'h1;
    T2[1166] = 2'h2;
    T2[1167] = 2'h2;
    T2[1168] = 2'h3;
    T2[1169] = 2'h0;
    T2[1170] = 2'h2;
    T2[1171] = 2'h2;
    T2[1172] = 2'h2;
    T2[1173] = 2'h3;
    T2[1174] = 2'h0;
    T2[1175] = 2'h3;
    T2[1176] = 2'h2;
    T2[1177] = 2'h2;
    T2[1178] = 2'h3;
    T2[1179] = 2'h0;
    T2[1180] = 2'h0;
    T2[1181] = 2'h3;
    T2[1182] = 2'h2;
    T2[1183] = 2'h3;
    T2[1184] = 2'h0;
    T2[1185] = 2'h1;
    T2[1186] = 2'h3;
    T2[1187] = 2'h2;
    T2[1188] = 2'h3;
    T2[1189] = 2'h0;
    T2[1190] = 2'h2;
    T2[1191] = 2'h3;
    T2[1192] = 2'h2;
    T2[1193] = 2'h3;
    T2[1194] = 2'h0;
    T2[1195] = 2'h3;
    T2[1196] = 2'h3;
    T2[1197] = 2'h2;
    T2[1198] = 2'h3;
    T2[1199] = 2'h0;
    T2[1200] = 2'h0;
    T2[1201] = 2'h0;
    T2[1202] = 2'h3;
    T2[1203] = 2'h3;
    T2[1204] = 2'h0;
    T2[1205] = 2'h1;
    T2[1206] = 2'h0;
    T2[1207] = 2'h3;
    T2[1208] = 2'h3;
    T2[1209] = 2'h0;
    T2[1210] = 2'h2;
    T2[1211] = 2'h0;
    T2[1212] = 2'h3;
    T2[1213] = 2'h3;
    T2[1214] = 2'h0;
    T2[1215] = 2'h3;
    T2[1216] = 2'h0;
    T2[1217] = 2'h3;
    T2[1218] = 2'h3;
    T2[1219] = 2'h0;
    T2[1220] = 2'h0;
    T2[1221] = 2'h1;
    T2[1222] = 2'h3;
    T2[1223] = 2'h3;
    T2[1224] = 2'h0;
    T2[1225] = 2'h1;
    T2[1226] = 2'h1;
    T2[1227] = 2'h3;
    T2[1228] = 2'h3;
    T2[1229] = 2'h0;
    T2[1230] = 2'h2;
    T2[1231] = 2'h1;
    T2[1232] = 2'h3;
    T2[1233] = 2'h3;
    T2[1234] = 2'h0;
    T2[1235] = 2'h3;
    T2[1236] = 2'h1;
    T2[1237] = 2'h3;
    T2[1238] = 2'h3;
    T2[1239] = 2'h0;
    T2[1240] = 2'h0;
    T2[1241] = 2'h2;
    T2[1242] = 2'h3;
    T2[1243] = 2'h3;
    T2[1244] = 2'h0;
    T2[1245] = 2'h1;
    T2[1246] = 2'h2;
    T2[1247] = 2'h3;
    T2[1248] = 2'h3;
    T2[1249] = 2'h0;
    T2[1250] = 2'h2;
    T2[1251] = 2'h2;
    T2[1252] = 2'h3;
    T2[1253] = 2'h3;
    T2[1254] = 2'h0;
    T2[1255] = 2'h3;
    T2[1256] = 2'h2;
    T2[1257] = 2'h3;
    T2[1258] = 2'h3;
    T2[1259] = 2'h0;
    T2[1260] = 2'h0;
    T2[1261] = 2'h3;
    T2[1262] = 2'h3;
    T2[1263] = 2'h3;
    T2[1264] = 2'h0;
    T2[1265] = 2'h1;
    T2[1266] = 2'h3;
    T2[1267] = 2'h3;
    T2[1268] = 2'h3;
    T2[1269] = 2'h0;
    T2[1270] = 2'h2;
    T2[1271] = 2'h3;
    T2[1272] = 2'h3;
    T2[1273] = 2'h3;
    T2[1274] = 2'h0;
    T2[1275] = 2'h3;
    T2[1276] = 2'h3;
    T2[1277] = 2'h3;
    T2[1278] = 2'h3;
    T2[1279] = 2'h0;
    T2[1280] = 2'h0;
    T2[1281] = 2'h0;
    T2[1282] = 2'h0;
    T2[1283] = 2'h0;
    T2[1284] = 2'h1;
    T2[1285] = 2'h1;
    T2[1286] = 2'h0;
    T2[1287] = 2'h0;
    T2[1288] = 2'h0;
    T2[1289] = 2'h1;
    T2[1290] = 2'h2;
    T2[1291] = 2'h0;
    T2[1292] = 2'h0;
    T2[1293] = 2'h0;
    T2[1294] = 2'h1;
    T2[1295] = 2'h3;
    T2[1296] = 2'h0;
    T2[1297] = 2'h0;
    T2[1298] = 2'h0;
    T2[1299] = 2'h1;
    T2[1300] = 2'h0;
    T2[1301] = 2'h1;
    T2[1302] = 2'h0;
    T2[1303] = 2'h0;
    T2[1304] = 2'h1;
    T2[1305] = 2'h1;
    T2[1306] = 2'h1;
    T2[1307] = 2'h0;
    T2[1308] = 2'h0;
    T2[1309] = 2'h1;
    T2[1310] = 2'h2;
    T2[1311] = 2'h1;
    T2[1312] = 2'h0;
    T2[1313] = 2'h0;
    T2[1314] = 2'h1;
    T2[1315] = 2'h3;
    T2[1316] = 2'h1;
    T2[1317] = 2'h0;
    T2[1318] = 2'h0;
    T2[1319] = 2'h1;
    T2[1320] = 2'h0;
    T2[1321] = 2'h2;
    T2[1322] = 2'h0;
    T2[1323] = 2'h0;
    T2[1324] = 2'h1;
    T2[1325] = 2'h1;
    T2[1326] = 2'h2;
    T2[1327] = 2'h0;
    T2[1328] = 2'h0;
    T2[1329] = 2'h1;
    T2[1330] = 2'h2;
    T2[1331] = 2'h2;
    T2[1332] = 2'h0;
    T2[1333] = 2'h0;
    T2[1334] = 2'h1;
    T2[1335] = 2'h3;
    T2[1336] = 2'h2;
    T2[1337] = 2'h0;
    T2[1338] = 2'h0;
    T2[1339] = 2'h1;
    T2[1340] = 2'h0;
    T2[1341] = 2'h3;
    T2[1342] = 2'h0;
    T2[1343] = 2'h0;
    T2[1344] = 2'h1;
    T2[1345] = 2'h1;
    T2[1346] = 2'h3;
    T2[1347] = 2'h0;
    T2[1348] = 2'h0;
    T2[1349] = 2'h1;
    T2[1350] = 2'h2;
    T2[1351] = 2'h3;
    T2[1352] = 2'h0;
    T2[1353] = 2'h0;
    T2[1354] = 2'h1;
    T2[1355] = 2'h3;
    T2[1356] = 2'h3;
    T2[1357] = 2'h0;
    T2[1358] = 2'h0;
    T2[1359] = 2'h1;
    T2[1360] = 2'h0;
    T2[1361] = 2'h0;
    T2[1362] = 2'h1;
    T2[1363] = 2'h0;
    T2[1364] = 2'h1;
    T2[1365] = 2'h1;
    T2[1366] = 2'h0;
    T2[1367] = 2'h1;
    T2[1368] = 2'h0;
    T2[1369] = 2'h1;
    T2[1370] = 2'h2;
    T2[1371] = 2'h0;
    T2[1372] = 2'h1;
    T2[1373] = 2'h0;
    T2[1374] = 2'h1;
    T2[1375] = 2'h3;
    T2[1376] = 2'h0;
    T2[1377] = 2'h1;
    T2[1378] = 2'h0;
    T2[1379] = 2'h1;
    T2[1380] = 2'h0;
    T2[1381] = 2'h1;
    T2[1382] = 2'h1;
    T2[1383] = 2'h0;
    T2[1384] = 2'h1;
    T2[1385] = 2'h1;
    T2[1386] = 2'h1;
    T2[1387] = 2'h1;
    T2[1388] = 2'h0;
    T2[1389] = 2'h1;
    T2[1390] = 2'h2;
    T2[1391] = 2'h1;
    T2[1392] = 2'h1;
    T2[1393] = 2'h0;
    T2[1394] = 2'h1;
    T2[1395] = 2'h3;
    T2[1396] = 2'h1;
    T2[1397] = 2'h1;
    T2[1398] = 2'h0;
    T2[1399] = 2'h1;
    T2[1400] = 2'h0;
    T2[1401] = 2'h2;
    T2[1402] = 2'h1;
    T2[1403] = 2'h0;
    T2[1404] = 2'h1;
    T2[1405] = 2'h1;
    T2[1406] = 2'h2;
    T2[1407] = 2'h1;
    T2[1408] = 2'h0;
    T2[1409] = 2'h1;
    T2[1410] = 2'h2;
    T2[1411] = 2'h2;
    T2[1412] = 2'h1;
    T2[1413] = 2'h0;
    T2[1414] = 2'h1;
    T2[1415] = 2'h3;
    T2[1416] = 2'h2;
    T2[1417] = 2'h1;
    T2[1418] = 2'h0;
    T2[1419] = 2'h1;
    T2[1420] = 2'h0;
    T2[1421] = 2'h3;
    T2[1422] = 2'h1;
    T2[1423] = 2'h0;
    T2[1424] = 2'h1;
    T2[1425] = 2'h1;
    T2[1426] = 2'h3;
    T2[1427] = 2'h1;
    T2[1428] = 2'h0;
    T2[1429] = 2'h1;
    T2[1430] = 2'h2;
    T2[1431] = 2'h3;
    T2[1432] = 2'h1;
    T2[1433] = 2'h0;
    T2[1434] = 2'h1;
    T2[1435] = 2'h3;
    T2[1436] = 2'h3;
    T2[1437] = 2'h1;
    T2[1438] = 2'h0;
    T2[1439] = 2'h1;
    T2[1440] = 2'h0;
    T2[1441] = 2'h0;
    T2[1442] = 2'h2;
    T2[1443] = 2'h0;
    T2[1444] = 2'h1;
    T2[1445] = 2'h1;
    T2[1446] = 2'h0;
    T2[1447] = 2'h2;
    T2[1448] = 2'h0;
    T2[1449] = 2'h1;
    T2[1450] = 2'h2;
    T2[1451] = 2'h0;
    T2[1452] = 2'h2;
    T2[1453] = 2'h0;
    T2[1454] = 2'h1;
    T2[1455] = 2'h3;
    T2[1456] = 2'h0;
    T2[1457] = 2'h2;
    T2[1458] = 2'h0;
    T2[1459] = 2'h1;
    T2[1460] = 2'h0;
    T2[1461] = 2'h1;
    T2[1462] = 2'h2;
    T2[1463] = 2'h0;
    T2[1464] = 2'h1;
    T2[1465] = 2'h1;
    T2[1466] = 2'h1;
    T2[1467] = 2'h2;
    T2[1468] = 2'h0;
    T2[1469] = 2'h1;
    T2[1470] = 2'h2;
    T2[1471] = 2'h1;
    T2[1472] = 2'h2;
    T2[1473] = 2'h0;
    T2[1474] = 2'h1;
    T2[1475] = 2'h3;
    T2[1476] = 2'h1;
    T2[1477] = 2'h2;
    T2[1478] = 2'h0;
    T2[1479] = 2'h1;
    T2[1480] = 2'h0;
    T2[1481] = 2'h2;
    T2[1482] = 2'h2;
    T2[1483] = 2'h0;
    T2[1484] = 2'h1;
    T2[1485] = 2'h1;
    T2[1486] = 2'h2;
    T2[1487] = 2'h2;
    T2[1488] = 2'h0;
    T2[1489] = 2'h1;
    T2[1490] = 2'h2;
    T2[1491] = 2'h2;
    T2[1492] = 2'h2;
    T2[1493] = 2'h0;
    T2[1494] = 2'h1;
    T2[1495] = 2'h3;
    T2[1496] = 2'h2;
    T2[1497] = 2'h2;
    T2[1498] = 2'h0;
    T2[1499] = 2'h1;
    T2[1500] = 2'h0;
    T2[1501] = 2'h3;
    T2[1502] = 2'h2;
    T2[1503] = 2'h0;
    T2[1504] = 2'h1;
    T2[1505] = 2'h1;
    T2[1506] = 2'h3;
    T2[1507] = 2'h2;
    T2[1508] = 2'h0;
    T2[1509] = 2'h1;
    T2[1510] = 2'h2;
    T2[1511] = 2'h3;
    T2[1512] = 2'h2;
    T2[1513] = 2'h0;
    T2[1514] = 2'h1;
    T2[1515] = 2'h3;
    T2[1516] = 2'h3;
    T2[1517] = 2'h2;
    T2[1518] = 2'h0;
    T2[1519] = 2'h1;
    T2[1520] = 2'h0;
    T2[1521] = 2'h0;
    T2[1522] = 2'h3;
    T2[1523] = 2'h0;
    T2[1524] = 2'h1;
    T2[1525] = 2'h1;
    T2[1526] = 2'h0;
    T2[1527] = 2'h3;
    T2[1528] = 2'h0;
    T2[1529] = 2'h1;
    T2[1530] = 2'h2;
    T2[1531] = 2'h0;
    T2[1532] = 2'h3;
    T2[1533] = 2'h0;
    T2[1534] = 2'h1;
    T2[1535] = 2'h3;
    T2[1536] = 2'h0;
    T2[1537] = 2'h3;
    T2[1538] = 2'h0;
    T2[1539] = 2'h1;
    T2[1540] = 2'h0;
    T2[1541] = 2'h1;
    T2[1542] = 2'h3;
    T2[1543] = 2'h0;
    T2[1544] = 2'h1;
    T2[1545] = 2'h1;
    T2[1546] = 2'h1;
    T2[1547] = 2'h3;
    T2[1548] = 2'h0;
    T2[1549] = 2'h1;
    T2[1550] = 2'h2;
    T2[1551] = 2'h1;
    T2[1552] = 2'h3;
    T2[1553] = 2'h0;
    T2[1554] = 2'h1;
    T2[1555] = 2'h3;
    T2[1556] = 2'h1;
    T2[1557] = 2'h3;
    T2[1558] = 2'h0;
    T2[1559] = 2'h1;
    T2[1560] = 2'h0;
    T2[1561] = 2'h2;
    T2[1562] = 2'h3;
    T2[1563] = 2'h0;
    T2[1564] = 2'h1;
    T2[1565] = 2'h1;
    T2[1566] = 2'h2;
    T2[1567] = 2'h3;
    T2[1568] = 2'h0;
    T2[1569] = 2'h1;
    T2[1570] = 2'h2;
    T2[1571] = 2'h2;
    T2[1572] = 2'h3;
    T2[1573] = 2'h0;
    T2[1574] = 2'h1;
    T2[1575] = 2'h3;
    T2[1576] = 2'h2;
    T2[1577] = 2'h3;
    T2[1578] = 2'h0;
    T2[1579] = 2'h1;
    T2[1580] = 2'h0;
    T2[1581] = 2'h3;
    T2[1582] = 2'h3;
    T2[1583] = 2'h0;
    T2[1584] = 2'h1;
    T2[1585] = 2'h1;
    T2[1586] = 2'h3;
    T2[1587] = 2'h3;
    T2[1588] = 2'h0;
    T2[1589] = 2'h1;
    T2[1590] = 2'h2;
    T2[1591] = 2'h3;
    T2[1592] = 2'h3;
    T2[1593] = 2'h0;
    T2[1594] = 2'h1;
    T2[1595] = 2'h3;
    T2[1596] = 2'h3;
    T2[1597] = 2'h3;
    T2[1598] = 2'h0;
    T2[1599] = 2'h1;
    T2[1600] = 2'h0;
    T2[1601] = 2'h0;
    T2[1602] = 2'h0;
    T2[1603] = 2'h1;
    T2[1604] = 2'h1;
    T2[1605] = 2'h1;
    T2[1606] = 2'h0;
    T2[1607] = 2'h0;
    T2[1608] = 2'h1;
    T2[1609] = 2'h1;
    T2[1610] = 2'h2;
    T2[1611] = 2'h0;
    T2[1612] = 2'h0;
    T2[1613] = 2'h1;
    T2[1614] = 2'h1;
    T2[1615] = 2'h3;
    T2[1616] = 2'h0;
    T2[1617] = 2'h0;
    T2[1618] = 2'h1;
    T2[1619] = 2'h1;
    T2[1620] = 2'h0;
    T2[1621] = 2'h1;
    T2[1622] = 2'h0;
    T2[1623] = 2'h1;
    T2[1624] = 2'h1;
    T2[1625] = 2'h1;
    T2[1626] = 2'h1;
    T2[1627] = 2'h0;
    T2[1628] = 2'h1;
    T2[1629] = 2'h1;
    T2[1630] = 2'h2;
    T2[1631] = 2'h1;
    T2[1632] = 2'h0;
    T2[1633] = 2'h1;
    T2[1634] = 2'h1;
    T2[1635] = 2'h3;
    T2[1636] = 2'h1;
    T2[1637] = 2'h0;
    T2[1638] = 2'h1;
    T2[1639] = 2'h1;
    T2[1640] = 2'h0;
    T2[1641] = 2'h2;
    T2[1642] = 2'h0;
    T2[1643] = 2'h1;
    T2[1644] = 2'h1;
    T2[1645] = 2'h1;
    T2[1646] = 2'h2;
    T2[1647] = 2'h0;
    T2[1648] = 2'h1;
    T2[1649] = 2'h1;
    T2[1650] = 2'h2;
    T2[1651] = 2'h2;
    T2[1652] = 2'h0;
    T2[1653] = 2'h1;
    T2[1654] = 2'h1;
    T2[1655] = 2'h3;
    T2[1656] = 2'h2;
    T2[1657] = 2'h0;
    T2[1658] = 2'h1;
    T2[1659] = 2'h1;
    T2[1660] = 2'h0;
    T2[1661] = 2'h3;
    T2[1662] = 2'h0;
    T2[1663] = 2'h1;
    T2[1664] = 2'h1;
    T2[1665] = 2'h1;
    T2[1666] = 2'h3;
    T2[1667] = 2'h0;
    T2[1668] = 2'h1;
    T2[1669] = 2'h1;
    T2[1670] = 2'h2;
    T2[1671] = 2'h3;
    T2[1672] = 2'h0;
    T2[1673] = 2'h1;
    T2[1674] = 2'h1;
    T2[1675] = 2'h3;
    T2[1676] = 2'h3;
    T2[1677] = 2'h0;
    T2[1678] = 2'h1;
    T2[1679] = 2'h1;
    T2[1680] = 2'h0;
    T2[1681] = 2'h0;
    T2[1682] = 2'h1;
    T2[1683] = 2'h1;
    T2[1684] = 2'h1;
    T2[1685] = 2'h1;
    T2[1686] = 2'h0;
    T2[1687] = 2'h1;
    T2[1688] = 2'h1;
    T2[1689] = 2'h1;
    T2[1690] = 2'h2;
    T2[1691] = 2'h0;
    T2[1692] = 2'h1;
    T2[1693] = 2'h1;
    T2[1694] = 2'h1;
    T2[1695] = 2'h3;
    T2[1696] = 2'h0;
    T2[1697] = 2'h1;
    T2[1698] = 2'h1;
    T2[1699] = 2'h1;
    T2[1700] = 2'h0;
    T2[1701] = 2'h1;
    T2[1702] = 2'h1;
    T2[1703] = 2'h1;
    T2[1704] = 2'h1;
    T2[1705] = 2'h1;
    T2[1706] = 2'h1;
    T2[1707] = 2'h1;
    T2[1708] = 2'h1;
    T2[1709] = 2'h1;
    T2[1710] = 2'h2;
    T2[1711] = 2'h1;
    T2[1712] = 2'h1;
    T2[1713] = 2'h1;
    T2[1714] = 2'h1;
    T2[1715] = 2'h3;
    T2[1716] = 2'h1;
    T2[1717] = 2'h1;
    T2[1718] = 2'h1;
    T2[1719] = 2'h1;
    T2[1720] = 2'h0;
    T2[1721] = 2'h2;
    T2[1722] = 2'h1;
    T2[1723] = 2'h1;
    T2[1724] = 2'h1;
    T2[1725] = 2'h1;
    T2[1726] = 2'h2;
    T2[1727] = 2'h1;
    T2[1728] = 2'h1;
    T2[1729] = 2'h1;
    T2[1730] = 2'h2;
    T2[1731] = 2'h2;
    T2[1732] = 2'h1;
    T2[1733] = 2'h1;
    T2[1734] = 2'h1;
    T2[1735] = 2'h3;
    T2[1736] = 2'h2;
    T2[1737] = 2'h1;
    T2[1738] = 2'h1;
    T2[1739] = 2'h1;
    T2[1740] = 2'h0;
    T2[1741] = 2'h3;
    T2[1742] = 2'h1;
    T2[1743] = 2'h1;
    T2[1744] = 2'h1;
    T2[1745] = 2'h1;
    T2[1746] = 2'h3;
    T2[1747] = 2'h1;
    T2[1748] = 2'h1;
    T2[1749] = 2'h1;
    T2[1750] = 2'h2;
    T2[1751] = 2'h3;
    T2[1752] = 2'h1;
    T2[1753] = 2'h1;
    T2[1754] = 2'h1;
    T2[1755] = 2'h3;
    T2[1756] = 2'h3;
    T2[1757] = 2'h1;
    T2[1758] = 2'h1;
    T2[1759] = 2'h1;
    T2[1760] = 2'h0;
    T2[1761] = 2'h0;
    T2[1762] = 2'h2;
    T2[1763] = 2'h1;
    T2[1764] = 2'h1;
    T2[1765] = 2'h1;
    T2[1766] = 2'h0;
    T2[1767] = 2'h2;
    T2[1768] = 2'h1;
    T2[1769] = 2'h1;
    T2[1770] = 2'h2;
    T2[1771] = 2'h0;
    T2[1772] = 2'h2;
    T2[1773] = 2'h1;
    T2[1774] = 2'h1;
    T2[1775] = 2'h3;
    T2[1776] = 2'h0;
    T2[1777] = 2'h2;
    T2[1778] = 2'h1;
    T2[1779] = 2'h1;
    T2[1780] = 2'h0;
    T2[1781] = 2'h1;
    T2[1782] = 2'h2;
    T2[1783] = 2'h1;
    T2[1784] = 2'h1;
    T2[1785] = 2'h1;
    T2[1786] = 2'h1;
    T2[1787] = 2'h2;
    T2[1788] = 2'h1;
    T2[1789] = 2'h1;
    T2[1790] = 2'h2;
    T2[1791] = 2'h1;
    T2[1792] = 2'h2;
    T2[1793] = 2'h1;
    T2[1794] = 2'h1;
    T2[1795] = 2'h3;
    T2[1796] = 2'h1;
    T2[1797] = 2'h2;
    T2[1798] = 2'h1;
    T2[1799] = 2'h1;
    T2[1800] = 2'h0;
    T2[1801] = 2'h2;
    T2[1802] = 2'h2;
    T2[1803] = 2'h1;
    T2[1804] = 2'h1;
    T2[1805] = 2'h1;
    T2[1806] = 2'h2;
    T2[1807] = 2'h2;
    T2[1808] = 2'h1;
    T2[1809] = 2'h1;
    T2[1810] = 2'h2;
    T2[1811] = 2'h2;
    T2[1812] = 2'h2;
    T2[1813] = 2'h1;
    T2[1814] = 2'h1;
    T2[1815] = 2'h3;
    T2[1816] = 2'h2;
    T2[1817] = 2'h2;
    T2[1818] = 2'h1;
    T2[1819] = 2'h1;
    T2[1820] = 2'h0;
    T2[1821] = 2'h3;
    T2[1822] = 2'h2;
    T2[1823] = 2'h1;
    T2[1824] = 2'h1;
    T2[1825] = 2'h1;
    T2[1826] = 2'h3;
    T2[1827] = 2'h2;
    T2[1828] = 2'h1;
    T2[1829] = 2'h1;
    T2[1830] = 2'h2;
    T2[1831] = 2'h3;
    T2[1832] = 2'h2;
    T2[1833] = 2'h1;
    T2[1834] = 2'h1;
    T2[1835] = 2'h3;
    T2[1836] = 2'h3;
    T2[1837] = 2'h2;
    T2[1838] = 2'h1;
    T2[1839] = 2'h1;
    T2[1840] = 2'h0;
    T2[1841] = 2'h0;
    T2[1842] = 2'h3;
    T2[1843] = 2'h1;
    T2[1844] = 2'h1;
    T2[1845] = 2'h1;
    T2[1846] = 2'h0;
    T2[1847] = 2'h3;
    T2[1848] = 2'h1;
    T2[1849] = 2'h1;
    T2[1850] = 2'h2;
    T2[1851] = 2'h0;
    T2[1852] = 2'h3;
    T2[1853] = 2'h1;
    T2[1854] = 2'h1;
    T2[1855] = 2'h3;
    T2[1856] = 2'h0;
    T2[1857] = 2'h3;
    T2[1858] = 2'h1;
    T2[1859] = 2'h1;
    T2[1860] = 2'h0;
    T2[1861] = 2'h1;
    T2[1862] = 2'h3;
    T2[1863] = 2'h1;
    T2[1864] = 2'h1;
    T2[1865] = 2'h1;
    T2[1866] = 2'h1;
    T2[1867] = 2'h3;
    T2[1868] = 2'h1;
    T2[1869] = 2'h1;
    T2[1870] = 2'h2;
    T2[1871] = 2'h1;
    T2[1872] = 2'h3;
    T2[1873] = 2'h1;
    T2[1874] = 2'h1;
    T2[1875] = 2'h3;
    T2[1876] = 2'h1;
    T2[1877] = 2'h3;
    T2[1878] = 2'h1;
    T2[1879] = 2'h1;
    T2[1880] = 2'h0;
    T2[1881] = 2'h2;
    T2[1882] = 2'h3;
    T2[1883] = 2'h1;
    T2[1884] = 2'h1;
    T2[1885] = 2'h1;
    T2[1886] = 2'h2;
    T2[1887] = 2'h3;
    T2[1888] = 2'h1;
    T2[1889] = 2'h1;
    T2[1890] = 2'h2;
    T2[1891] = 2'h2;
    T2[1892] = 2'h3;
    T2[1893] = 2'h1;
    T2[1894] = 2'h1;
    T2[1895] = 2'h3;
    T2[1896] = 2'h2;
    T2[1897] = 2'h3;
    T2[1898] = 2'h1;
    T2[1899] = 2'h1;
    T2[1900] = 2'h0;
    T2[1901] = 2'h3;
    T2[1902] = 2'h3;
    T2[1903] = 2'h1;
    T2[1904] = 2'h1;
    T2[1905] = 2'h1;
    T2[1906] = 2'h3;
    T2[1907] = 2'h3;
    T2[1908] = 2'h1;
    T2[1909] = 2'h1;
    T2[1910] = 2'h2;
    T2[1911] = 2'h3;
    T2[1912] = 2'h3;
    T2[1913] = 2'h1;
    T2[1914] = 2'h1;
    T2[1915] = 2'h3;
    T2[1916] = 2'h3;
    T2[1917] = 2'h3;
    T2[1918] = 2'h1;
    T2[1919] = 2'h1;
    T2[1920] = 2'h0;
    T2[1921] = 2'h0;
    T2[1922] = 2'h0;
    T2[1923] = 2'h2;
    T2[1924] = 2'h1;
    T2[1925] = 2'h1;
    T2[1926] = 2'h0;
    T2[1927] = 2'h0;
    T2[1928] = 2'h2;
    T2[1929] = 2'h1;
    T2[1930] = 2'h2;
    T2[1931] = 2'h0;
    T2[1932] = 2'h0;
    T2[1933] = 2'h2;
    T2[1934] = 2'h1;
    T2[1935] = 2'h3;
    T2[1936] = 2'h0;
    T2[1937] = 2'h0;
    T2[1938] = 2'h2;
    T2[1939] = 2'h1;
    T2[1940] = 2'h0;
    T2[1941] = 2'h1;
    T2[1942] = 2'h0;
    T2[1943] = 2'h2;
    T2[1944] = 2'h1;
    T2[1945] = 2'h1;
    T2[1946] = 2'h1;
    T2[1947] = 2'h0;
    T2[1948] = 2'h2;
    T2[1949] = 2'h1;
    T2[1950] = 2'h2;
    T2[1951] = 2'h1;
    T2[1952] = 2'h0;
    T2[1953] = 2'h2;
    T2[1954] = 2'h1;
    T2[1955] = 2'h3;
    T2[1956] = 2'h1;
    T2[1957] = 2'h0;
    T2[1958] = 2'h2;
    T2[1959] = 2'h1;
    T2[1960] = 2'h0;
    T2[1961] = 2'h2;
    T2[1962] = 2'h0;
    T2[1963] = 2'h2;
    T2[1964] = 2'h1;
    T2[1965] = 2'h1;
    T2[1966] = 2'h2;
    T2[1967] = 2'h0;
    T2[1968] = 2'h2;
    T2[1969] = 2'h1;
    T2[1970] = 2'h2;
    T2[1971] = 2'h2;
    T2[1972] = 2'h0;
    T2[1973] = 2'h2;
    T2[1974] = 2'h1;
    T2[1975] = 2'h3;
    T2[1976] = 2'h2;
    T2[1977] = 2'h0;
    T2[1978] = 2'h2;
    T2[1979] = 2'h1;
    T2[1980] = 2'h0;
    T2[1981] = 2'h3;
    T2[1982] = 2'h0;
    T2[1983] = 2'h2;
    T2[1984] = 2'h1;
    T2[1985] = 2'h1;
    T2[1986] = 2'h3;
    T2[1987] = 2'h0;
    T2[1988] = 2'h2;
    T2[1989] = 2'h1;
    T2[1990] = 2'h2;
    T2[1991] = 2'h3;
    T2[1992] = 2'h0;
    T2[1993] = 2'h2;
    T2[1994] = 2'h1;
    T2[1995] = 2'h3;
    T2[1996] = 2'h3;
    T2[1997] = 2'h0;
    T2[1998] = 2'h2;
    T2[1999] = 2'h1;
    T2[2000] = 2'h0;
    T2[2001] = 2'h0;
    T2[2002] = 2'h1;
    T2[2003] = 2'h2;
    T2[2004] = 2'h1;
    T2[2005] = 2'h1;
    T2[2006] = 2'h0;
    T2[2007] = 2'h1;
    T2[2008] = 2'h2;
    T2[2009] = 2'h1;
    T2[2010] = 2'h2;
    T2[2011] = 2'h0;
    T2[2012] = 2'h1;
    T2[2013] = 2'h2;
    T2[2014] = 2'h1;
    T2[2015] = 2'h3;
    T2[2016] = 2'h0;
    T2[2017] = 2'h1;
    T2[2018] = 2'h2;
    T2[2019] = 2'h1;
    T2[2020] = 2'h0;
    T2[2021] = 2'h1;
    T2[2022] = 2'h1;
    T2[2023] = 2'h2;
    T2[2024] = 2'h1;
    T2[2025] = 2'h1;
    T2[2026] = 2'h1;
    T2[2027] = 2'h1;
    T2[2028] = 2'h2;
    T2[2029] = 2'h1;
    T2[2030] = 2'h2;
    T2[2031] = 2'h1;
    T2[2032] = 2'h1;
    T2[2033] = 2'h2;
    T2[2034] = 2'h1;
    T2[2035] = 2'h3;
    T2[2036] = 2'h1;
    T2[2037] = 2'h1;
    T2[2038] = 2'h2;
    T2[2039] = 2'h1;
    T2[2040] = 2'h0;
    T2[2041] = 2'h2;
    T2[2042] = 2'h1;
    T2[2043] = 2'h2;
    T2[2044] = 2'h1;
    T2[2045] = 2'h1;
    T2[2046] = 2'h2;
    T2[2047] = 2'h1;
    T2[2048] = 2'h2;
    T2[2049] = 2'h1;
    T2[2050] = 2'h2;
    T2[2051] = 2'h2;
    T2[2052] = 2'h1;
    T2[2053] = 2'h2;
    T2[2054] = 2'h1;
    T2[2055] = 2'h3;
    T2[2056] = 2'h2;
    T2[2057] = 2'h1;
    T2[2058] = 2'h2;
    T2[2059] = 2'h1;
    T2[2060] = 2'h0;
    T2[2061] = 2'h3;
    T2[2062] = 2'h1;
    T2[2063] = 2'h2;
    T2[2064] = 2'h1;
    T2[2065] = 2'h1;
    T2[2066] = 2'h3;
    T2[2067] = 2'h1;
    T2[2068] = 2'h2;
    T2[2069] = 2'h1;
    T2[2070] = 2'h2;
    T2[2071] = 2'h3;
    T2[2072] = 2'h1;
    T2[2073] = 2'h2;
    T2[2074] = 2'h1;
    T2[2075] = 2'h3;
    T2[2076] = 2'h3;
    T2[2077] = 2'h1;
    T2[2078] = 2'h2;
    T2[2079] = 2'h1;
    T2[2080] = 2'h0;
    T2[2081] = 2'h0;
    T2[2082] = 2'h2;
    T2[2083] = 2'h2;
    T2[2084] = 2'h1;
    T2[2085] = 2'h1;
    T2[2086] = 2'h0;
    T2[2087] = 2'h2;
    T2[2088] = 2'h2;
    T2[2089] = 2'h1;
    T2[2090] = 2'h2;
    T2[2091] = 2'h0;
    T2[2092] = 2'h2;
    T2[2093] = 2'h2;
    T2[2094] = 2'h1;
    T2[2095] = 2'h3;
    T2[2096] = 2'h0;
    T2[2097] = 2'h2;
    T2[2098] = 2'h2;
    T2[2099] = 2'h1;
    T2[2100] = 2'h0;
    T2[2101] = 2'h1;
    T2[2102] = 2'h2;
    T2[2103] = 2'h2;
    T2[2104] = 2'h1;
    T2[2105] = 2'h1;
    T2[2106] = 2'h1;
    T2[2107] = 2'h2;
    T2[2108] = 2'h2;
    T2[2109] = 2'h1;
    T2[2110] = 2'h2;
    T2[2111] = 2'h1;
    T2[2112] = 2'h2;
    T2[2113] = 2'h2;
    T2[2114] = 2'h1;
    T2[2115] = 2'h3;
    T2[2116] = 2'h1;
    T2[2117] = 2'h2;
    T2[2118] = 2'h2;
    T2[2119] = 2'h1;
    T2[2120] = 2'h0;
    T2[2121] = 2'h2;
    T2[2122] = 2'h2;
    T2[2123] = 2'h2;
    T2[2124] = 2'h1;
    T2[2125] = 2'h1;
    T2[2126] = 2'h2;
    T2[2127] = 2'h2;
    T2[2128] = 2'h2;
    T2[2129] = 2'h1;
    T2[2130] = 2'h2;
    T2[2131] = 2'h2;
    T2[2132] = 2'h2;
    T2[2133] = 2'h2;
    T2[2134] = 2'h1;
    T2[2135] = 2'h3;
    T2[2136] = 2'h2;
    T2[2137] = 2'h2;
    T2[2138] = 2'h2;
    T2[2139] = 2'h1;
    T2[2140] = 2'h0;
    T2[2141] = 2'h3;
    T2[2142] = 2'h2;
    T2[2143] = 2'h2;
    T2[2144] = 2'h1;
    T2[2145] = 2'h1;
    T2[2146] = 2'h3;
    T2[2147] = 2'h2;
    T2[2148] = 2'h2;
    T2[2149] = 2'h1;
    T2[2150] = 2'h2;
    T2[2151] = 2'h3;
    T2[2152] = 2'h2;
    T2[2153] = 2'h2;
    T2[2154] = 2'h1;
    T2[2155] = 2'h3;
    T2[2156] = 2'h3;
    T2[2157] = 2'h2;
    T2[2158] = 2'h2;
    T2[2159] = 2'h1;
    T2[2160] = 2'h0;
    T2[2161] = 2'h0;
    T2[2162] = 2'h3;
    T2[2163] = 2'h2;
    T2[2164] = 2'h1;
    T2[2165] = 2'h1;
    T2[2166] = 2'h0;
    T2[2167] = 2'h3;
    T2[2168] = 2'h2;
    T2[2169] = 2'h1;
    T2[2170] = 2'h2;
    T2[2171] = 2'h0;
    T2[2172] = 2'h3;
    T2[2173] = 2'h2;
    T2[2174] = 2'h1;
    T2[2175] = 2'h3;
    T2[2176] = 2'h0;
    T2[2177] = 2'h3;
    T2[2178] = 2'h2;
    T2[2179] = 2'h1;
    T2[2180] = 2'h0;
    T2[2181] = 2'h1;
    T2[2182] = 2'h3;
    T2[2183] = 2'h2;
    T2[2184] = 2'h1;
    T2[2185] = 2'h1;
    T2[2186] = 2'h1;
    T2[2187] = 2'h3;
    T2[2188] = 2'h2;
    T2[2189] = 2'h1;
    T2[2190] = 2'h2;
    T2[2191] = 2'h1;
    T2[2192] = 2'h3;
    T2[2193] = 2'h2;
    T2[2194] = 2'h1;
    T2[2195] = 2'h3;
    T2[2196] = 2'h1;
    T2[2197] = 2'h3;
    T2[2198] = 2'h2;
    T2[2199] = 2'h1;
    T2[2200] = 2'h0;
    T2[2201] = 2'h2;
    T2[2202] = 2'h3;
    T2[2203] = 2'h2;
    T2[2204] = 2'h1;
    T2[2205] = 2'h1;
    T2[2206] = 2'h2;
    T2[2207] = 2'h3;
    T2[2208] = 2'h2;
    T2[2209] = 2'h1;
    T2[2210] = 2'h2;
    T2[2211] = 2'h2;
    T2[2212] = 2'h3;
    T2[2213] = 2'h2;
    T2[2214] = 2'h1;
    T2[2215] = 2'h3;
    T2[2216] = 2'h2;
    T2[2217] = 2'h3;
    T2[2218] = 2'h2;
    T2[2219] = 2'h1;
    T2[2220] = 2'h0;
    T2[2221] = 2'h3;
    T2[2222] = 2'h3;
    T2[2223] = 2'h2;
    T2[2224] = 2'h1;
    T2[2225] = 2'h1;
    T2[2226] = 2'h3;
    T2[2227] = 2'h3;
    T2[2228] = 2'h2;
    T2[2229] = 2'h1;
    T2[2230] = 2'h2;
    T2[2231] = 2'h3;
    T2[2232] = 2'h3;
    T2[2233] = 2'h2;
    T2[2234] = 2'h1;
    T2[2235] = 2'h3;
    T2[2236] = 2'h3;
    T2[2237] = 2'h3;
    T2[2238] = 2'h2;
    T2[2239] = 2'h1;
    T2[2240] = 2'h0;
    T2[2241] = 2'h0;
    T2[2242] = 2'h0;
    T2[2243] = 2'h3;
    T2[2244] = 2'h1;
    T2[2245] = 2'h1;
    T2[2246] = 2'h0;
    T2[2247] = 2'h0;
    T2[2248] = 2'h3;
    T2[2249] = 2'h1;
    T2[2250] = 2'h2;
    T2[2251] = 2'h0;
    T2[2252] = 2'h0;
    T2[2253] = 2'h3;
    T2[2254] = 2'h1;
    T2[2255] = 2'h3;
    T2[2256] = 2'h0;
    T2[2257] = 2'h0;
    T2[2258] = 2'h3;
    T2[2259] = 2'h1;
    T2[2260] = 2'h0;
    T2[2261] = 2'h1;
    T2[2262] = 2'h0;
    T2[2263] = 2'h3;
    T2[2264] = 2'h1;
    T2[2265] = 2'h1;
    T2[2266] = 2'h1;
    T2[2267] = 2'h0;
    T2[2268] = 2'h3;
    T2[2269] = 2'h1;
    T2[2270] = 2'h2;
    T2[2271] = 2'h1;
    T2[2272] = 2'h0;
    T2[2273] = 2'h3;
    T2[2274] = 2'h1;
    T2[2275] = 2'h3;
    T2[2276] = 2'h1;
    T2[2277] = 2'h0;
    T2[2278] = 2'h3;
    T2[2279] = 2'h1;
    T2[2280] = 2'h0;
    T2[2281] = 2'h2;
    T2[2282] = 2'h0;
    T2[2283] = 2'h3;
    T2[2284] = 2'h1;
    T2[2285] = 2'h1;
    T2[2286] = 2'h2;
    T2[2287] = 2'h0;
    T2[2288] = 2'h3;
    T2[2289] = 2'h1;
    T2[2290] = 2'h2;
    T2[2291] = 2'h2;
    T2[2292] = 2'h0;
    T2[2293] = 2'h3;
    T2[2294] = 2'h1;
    T2[2295] = 2'h3;
    T2[2296] = 2'h2;
    T2[2297] = 2'h0;
    T2[2298] = 2'h3;
    T2[2299] = 2'h1;
    T2[2300] = 2'h0;
    T2[2301] = 2'h3;
    T2[2302] = 2'h0;
    T2[2303] = 2'h3;
    T2[2304] = 2'h1;
    T2[2305] = 2'h1;
    T2[2306] = 2'h3;
    T2[2307] = 2'h0;
    T2[2308] = 2'h3;
    T2[2309] = 2'h1;
    T2[2310] = 2'h2;
    T2[2311] = 2'h3;
    T2[2312] = 2'h0;
    T2[2313] = 2'h3;
    T2[2314] = 2'h1;
    T2[2315] = 2'h3;
    T2[2316] = 2'h3;
    T2[2317] = 2'h0;
    T2[2318] = 2'h3;
    T2[2319] = 2'h1;
    T2[2320] = 2'h0;
    T2[2321] = 2'h0;
    T2[2322] = 2'h1;
    T2[2323] = 2'h3;
    T2[2324] = 2'h1;
    T2[2325] = 2'h1;
    T2[2326] = 2'h0;
    T2[2327] = 2'h1;
    T2[2328] = 2'h3;
    T2[2329] = 2'h1;
    T2[2330] = 2'h2;
    T2[2331] = 2'h0;
    T2[2332] = 2'h1;
    T2[2333] = 2'h3;
    T2[2334] = 2'h1;
    T2[2335] = 2'h3;
    T2[2336] = 2'h0;
    T2[2337] = 2'h1;
    T2[2338] = 2'h3;
    T2[2339] = 2'h1;
    T2[2340] = 2'h0;
    T2[2341] = 2'h1;
    T2[2342] = 2'h1;
    T2[2343] = 2'h3;
    T2[2344] = 2'h1;
    T2[2345] = 2'h1;
    T2[2346] = 2'h1;
    T2[2347] = 2'h1;
    T2[2348] = 2'h3;
    T2[2349] = 2'h1;
    T2[2350] = 2'h2;
    T2[2351] = 2'h1;
    T2[2352] = 2'h1;
    T2[2353] = 2'h3;
    T2[2354] = 2'h1;
    T2[2355] = 2'h3;
    T2[2356] = 2'h1;
    T2[2357] = 2'h1;
    T2[2358] = 2'h3;
    T2[2359] = 2'h1;
    T2[2360] = 2'h0;
    T2[2361] = 2'h2;
    T2[2362] = 2'h1;
    T2[2363] = 2'h3;
    T2[2364] = 2'h1;
    T2[2365] = 2'h1;
    T2[2366] = 2'h2;
    T2[2367] = 2'h1;
    T2[2368] = 2'h3;
    T2[2369] = 2'h1;
    T2[2370] = 2'h2;
    T2[2371] = 2'h2;
    T2[2372] = 2'h1;
    T2[2373] = 2'h3;
    T2[2374] = 2'h1;
    T2[2375] = 2'h3;
    T2[2376] = 2'h2;
    T2[2377] = 2'h1;
    T2[2378] = 2'h3;
    T2[2379] = 2'h1;
    T2[2380] = 2'h0;
    T2[2381] = 2'h3;
    T2[2382] = 2'h1;
    T2[2383] = 2'h3;
    T2[2384] = 2'h1;
    T2[2385] = 2'h1;
    T2[2386] = 2'h3;
    T2[2387] = 2'h1;
    T2[2388] = 2'h3;
    T2[2389] = 2'h1;
    T2[2390] = 2'h2;
    T2[2391] = 2'h3;
    T2[2392] = 2'h1;
    T2[2393] = 2'h3;
    T2[2394] = 2'h1;
    T2[2395] = 2'h3;
    T2[2396] = 2'h3;
    T2[2397] = 2'h1;
    T2[2398] = 2'h3;
    T2[2399] = 2'h1;
    T2[2400] = 2'h0;
    T2[2401] = 2'h0;
    T2[2402] = 2'h2;
    T2[2403] = 2'h3;
    T2[2404] = 2'h1;
    T2[2405] = 2'h1;
    T2[2406] = 2'h0;
    T2[2407] = 2'h2;
    T2[2408] = 2'h3;
    T2[2409] = 2'h1;
    T2[2410] = 2'h2;
    T2[2411] = 2'h0;
    T2[2412] = 2'h2;
    T2[2413] = 2'h3;
    T2[2414] = 2'h1;
    T2[2415] = 2'h3;
    T2[2416] = 2'h0;
    T2[2417] = 2'h2;
    T2[2418] = 2'h3;
    T2[2419] = 2'h1;
    T2[2420] = 2'h0;
    T2[2421] = 2'h1;
    T2[2422] = 2'h2;
    T2[2423] = 2'h3;
    T2[2424] = 2'h1;
    T2[2425] = 2'h1;
    T2[2426] = 2'h1;
    T2[2427] = 2'h2;
    T2[2428] = 2'h3;
    T2[2429] = 2'h1;
    T2[2430] = 2'h2;
    T2[2431] = 2'h1;
    T2[2432] = 2'h2;
    T2[2433] = 2'h3;
    T2[2434] = 2'h1;
    T2[2435] = 2'h3;
    T2[2436] = 2'h1;
    T2[2437] = 2'h2;
    T2[2438] = 2'h3;
    T2[2439] = 2'h1;
    T2[2440] = 2'h0;
    T2[2441] = 2'h2;
    T2[2442] = 2'h2;
    T2[2443] = 2'h3;
    T2[2444] = 2'h1;
    T2[2445] = 2'h1;
    T2[2446] = 2'h2;
    T2[2447] = 2'h2;
    T2[2448] = 2'h3;
    T2[2449] = 2'h1;
    T2[2450] = 2'h2;
    T2[2451] = 2'h2;
    T2[2452] = 2'h2;
    T2[2453] = 2'h3;
    T2[2454] = 2'h1;
    T2[2455] = 2'h3;
    T2[2456] = 2'h2;
    T2[2457] = 2'h2;
    T2[2458] = 2'h3;
    T2[2459] = 2'h1;
    T2[2460] = 2'h0;
    T2[2461] = 2'h3;
    T2[2462] = 2'h2;
    T2[2463] = 2'h3;
    T2[2464] = 2'h1;
    T2[2465] = 2'h1;
    T2[2466] = 2'h3;
    T2[2467] = 2'h2;
    T2[2468] = 2'h3;
    T2[2469] = 2'h1;
    T2[2470] = 2'h2;
    T2[2471] = 2'h3;
    T2[2472] = 2'h2;
    T2[2473] = 2'h3;
    T2[2474] = 2'h1;
    T2[2475] = 2'h3;
    T2[2476] = 2'h3;
    T2[2477] = 2'h2;
    T2[2478] = 2'h3;
    T2[2479] = 2'h1;
    T2[2480] = 2'h0;
    T2[2481] = 2'h0;
    T2[2482] = 2'h3;
    T2[2483] = 2'h3;
    T2[2484] = 2'h1;
    T2[2485] = 2'h1;
    T2[2486] = 2'h0;
    T2[2487] = 2'h3;
    T2[2488] = 2'h3;
    T2[2489] = 2'h1;
    T2[2490] = 2'h2;
    T2[2491] = 2'h0;
    T2[2492] = 2'h3;
    T2[2493] = 2'h3;
    T2[2494] = 2'h1;
    T2[2495] = 2'h3;
    T2[2496] = 2'h0;
    T2[2497] = 2'h3;
    T2[2498] = 2'h3;
    T2[2499] = 2'h1;
    T2[2500] = 2'h0;
    T2[2501] = 2'h1;
    T2[2502] = 2'h3;
    T2[2503] = 2'h3;
    T2[2504] = 2'h1;
    T2[2505] = 2'h1;
    T2[2506] = 2'h1;
    T2[2507] = 2'h3;
    T2[2508] = 2'h3;
    T2[2509] = 2'h1;
    T2[2510] = 2'h2;
    T2[2511] = 2'h1;
    T2[2512] = 2'h3;
    T2[2513] = 2'h3;
    T2[2514] = 2'h1;
    T2[2515] = 2'h3;
    T2[2516] = 2'h1;
    T2[2517] = 2'h3;
    T2[2518] = 2'h3;
    T2[2519] = 2'h1;
    T2[2520] = 2'h0;
    T2[2521] = 2'h2;
    T2[2522] = 2'h3;
    T2[2523] = 2'h3;
    T2[2524] = 2'h1;
    T2[2525] = 2'h1;
    T2[2526] = 2'h2;
    T2[2527] = 2'h3;
    T2[2528] = 2'h3;
    T2[2529] = 2'h1;
    T2[2530] = 2'h2;
    T2[2531] = 2'h2;
    T2[2532] = 2'h3;
    T2[2533] = 2'h3;
    T2[2534] = 2'h1;
    T2[2535] = 2'h3;
    T2[2536] = 2'h2;
    T2[2537] = 2'h3;
    T2[2538] = 2'h3;
    T2[2539] = 2'h1;
    T2[2540] = 2'h0;
    T2[2541] = 2'h3;
    T2[2542] = 2'h3;
    T2[2543] = 2'h3;
    T2[2544] = 2'h1;
    T2[2545] = 2'h1;
    T2[2546] = 2'h3;
    T2[2547] = 2'h3;
    T2[2548] = 2'h3;
    T2[2549] = 2'h1;
    T2[2550] = 2'h2;
    T2[2551] = 2'h3;
    T2[2552] = 2'h3;
    T2[2553] = 2'h3;
    T2[2554] = 2'h1;
    T2[2555] = 2'h3;
    T2[2556] = 2'h3;
    T2[2557] = 2'h3;
    T2[2558] = 2'h3;
    T2[2559] = 2'h1;
    T2[2560] = 2'h0;
    T2[2561] = 2'h0;
    T2[2562] = 2'h0;
    T2[2563] = 2'h0;
    T2[2564] = 2'h2;
    T2[2565] = 2'h1;
    T2[2566] = 2'h0;
    T2[2567] = 2'h0;
    T2[2568] = 2'h0;
    T2[2569] = 2'h2;
    T2[2570] = 2'h2;
    T2[2571] = 2'h0;
    T2[2572] = 2'h0;
    T2[2573] = 2'h0;
    T2[2574] = 2'h2;
    T2[2575] = 2'h3;
    T2[2576] = 2'h0;
    T2[2577] = 2'h0;
    T2[2578] = 2'h0;
    T2[2579] = 2'h2;
    T2[2580] = 2'h0;
    T2[2581] = 2'h1;
    T2[2582] = 2'h0;
    T2[2583] = 2'h0;
    T2[2584] = 2'h2;
    T2[2585] = 2'h1;
    T2[2586] = 2'h1;
    T2[2587] = 2'h0;
    T2[2588] = 2'h0;
    T2[2589] = 2'h2;
    T2[2590] = 2'h2;
    T2[2591] = 2'h1;
    T2[2592] = 2'h0;
    T2[2593] = 2'h0;
    T2[2594] = 2'h2;
    T2[2595] = 2'h3;
    T2[2596] = 2'h1;
    T2[2597] = 2'h0;
    T2[2598] = 2'h0;
    T2[2599] = 2'h2;
    T2[2600] = 2'h0;
    T2[2601] = 2'h2;
    T2[2602] = 2'h0;
    T2[2603] = 2'h0;
    T2[2604] = 2'h2;
    T2[2605] = 2'h1;
    T2[2606] = 2'h2;
    T2[2607] = 2'h0;
    T2[2608] = 2'h0;
    T2[2609] = 2'h2;
    T2[2610] = 2'h2;
    T2[2611] = 2'h2;
    T2[2612] = 2'h0;
    T2[2613] = 2'h0;
    T2[2614] = 2'h2;
    T2[2615] = 2'h3;
    T2[2616] = 2'h2;
    T2[2617] = 2'h0;
    T2[2618] = 2'h0;
    T2[2619] = 2'h2;
    T2[2620] = 2'h0;
    T2[2621] = 2'h3;
    T2[2622] = 2'h0;
    T2[2623] = 2'h0;
    T2[2624] = 2'h2;
    T2[2625] = 2'h1;
    T2[2626] = 2'h3;
    T2[2627] = 2'h0;
    T2[2628] = 2'h0;
    T2[2629] = 2'h2;
    T2[2630] = 2'h2;
    T2[2631] = 2'h3;
    T2[2632] = 2'h0;
    T2[2633] = 2'h0;
    T2[2634] = 2'h2;
    T2[2635] = 2'h3;
    T2[2636] = 2'h3;
    T2[2637] = 2'h0;
    T2[2638] = 2'h0;
    T2[2639] = 2'h2;
    T2[2640] = 2'h0;
    T2[2641] = 2'h0;
    T2[2642] = 2'h1;
    T2[2643] = 2'h0;
    T2[2644] = 2'h2;
    T2[2645] = 2'h1;
    T2[2646] = 2'h0;
    T2[2647] = 2'h1;
    T2[2648] = 2'h0;
    T2[2649] = 2'h2;
    T2[2650] = 2'h2;
    T2[2651] = 2'h0;
    T2[2652] = 2'h1;
    T2[2653] = 2'h0;
    T2[2654] = 2'h2;
    T2[2655] = 2'h3;
    T2[2656] = 2'h0;
    T2[2657] = 2'h1;
    T2[2658] = 2'h0;
    T2[2659] = 2'h2;
    T2[2660] = 2'h0;
    T2[2661] = 2'h1;
    T2[2662] = 2'h1;
    T2[2663] = 2'h0;
    T2[2664] = 2'h2;
    T2[2665] = 2'h1;
    T2[2666] = 2'h1;
    T2[2667] = 2'h1;
    T2[2668] = 2'h0;
    T2[2669] = 2'h2;
    T2[2670] = 2'h2;
    T2[2671] = 2'h1;
    T2[2672] = 2'h1;
    T2[2673] = 2'h0;
    T2[2674] = 2'h2;
    T2[2675] = 2'h3;
    T2[2676] = 2'h1;
    T2[2677] = 2'h1;
    T2[2678] = 2'h0;
    T2[2679] = 2'h2;
    T2[2680] = 2'h0;
    T2[2681] = 2'h2;
    T2[2682] = 2'h1;
    T2[2683] = 2'h0;
    T2[2684] = 2'h2;
    T2[2685] = 2'h1;
    T2[2686] = 2'h2;
    T2[2687] = 2'h1;
    T2[2688] = 2'h0;
    T2[2689] = 2'h2;
    T2[2690] = 2'h2;
    T2[2691] = 2'h2;
    T2[2692] = 2'h1;
    T2[2693] = 2'h0;
    T2[2694] = 2'h2;
    T2[2695] = 2'h3;
    T2[2696] = 2'h2;
    T2[2697] = 2'h1;
    T2[2698] = 2'h0;
    T2[2699] = 2'h2;
    T2[2700] = 2'h0;
    T2[2701] = 2'h3;
    T2[2702] = 2'h1;
    T2[2703] = 2'h0;
    T2[2704] = 2'h2;
    T2[2705] = 2'h1;
    T2[2706] = 2'h3;
    T2[2707] = 2'h1;
    T2[2708] = 2'h0;
    T2[2709] = 2'h2;
    T2[2710] = 2'h2;
    T2[2711] = 2'h3;
    T2[2712] = 2'h1;
    T2[2713] = 2'h0;
    T2[2714] = 2'h2;
    T2[2715] = 2'h3;
    T2[2716] = 2'h3;
    T2[2717] = 2'h1;
    T2[2718] = 2'h0;
    T2[2719] = 2'h2;
    T2[2720] = 2'h0;
    T2[2721] = 2'h0;
    T2[2722] = 2'h2;
    T2[2723] = 2'h0;
    T2[2724] = 2'h2;
    T2[2725] = 2'h1;
    T2[2726] = 2'h0;
    T2[2727] = 2'h2;
    T2[2728] = 2'h0;
    T2[2729] = 2'h2;
    T2[2730] = 2'h2;
    T2[2731] = 2'h0;
    T2[2732] = 2'h2;
    T2[2733] = 2'h0;
    T2[2734] = 2'h2;
    T2[2735] = 2'h3;
    T2[2736] = 2'h0;
    T2[2737] = 2'h2;
    T2[2738] = 2'h0;
    T2[2739] = 2'h2;
    T2[2740] = 2'h0;
    T2[2741] = 2'h1;
    T2[2742] = 2'h2;
    T2[2743] = 2'h0;
    T2[2744] = 2'h2;
    T2[2745] = 2'h1;
    T2[2746] = 2'h1;
    T2[2747] = 2'h2;
    T2[2748] = 2'h0;
    T2[2749] = 2'h2;
    T2[2750] = 2'h2;
    T2[2751] = 2'h1;
    T2[2752] = 2'h2;
    T2[2753] = 2'h0;
    T2[2754] = 2'h2;
    T2[2755] = 2'h3;
    T2[2756] = 2'h1;
    T2[2757] = 2'h2;
    T2[2758] = 2'h0;
    T2[2759] = 2'h2;
    T2[2760] = 2'h0;
    T2[2761] = 2'h2;
    T2[2762] = 2'h2;
    T2[2763] = 2'h0;
    T2[2764] = 2'h2;
    T2[2765] = 2'h1;
    T2[2766] = 2'h2;
    T2[2767] = 2'h2;
    T2[2768] = 2'h0;
    T2[2769] = 2'h2;
    T2[2770] = 2'h2;
    T2[2771] = 2'h2;
    T2[2772] = 2'h2;
    T2[2773] = 2'h0;
    T2[2774] = 2'h2;
    T2[2775] = 2'h3;
    T2[2776] = 2'h2;
    T2[2777] = 2'h2;
    T2[2778] = 2'h0;
    T2[2779] = 2'h2;
    T2[2780] = 2'h0;
    T2[2781] = 2'h3;
    T2[2782] = 2'h2;
    T2[2783] = 2'h0;
    T2[2784] = 2'h2;
    T2[2785] = 2'h1;
    T2[2786] = 2'h3;
    T2[2787] = 2'h2;
    T2[2788] = 2'h0;
    T2[2789] = 2'h2;
    T2[2790] = 2'h2;
    T2[2791] = 2'h3;
    T2[2792] = 2'h2;
    T2[2793] = 2'h0;
    T2[2794] = 2'h2;
    T2[2795] = 2'h3;
    T2[2796] = 2'h3;
    T2[2797] = 2'h2;
    T2[2798] = 2'h0;
    T2[2799] = 2'h2;
    T2[2800] = 2'h0;
    T2[2801] = 2'h0;
    T2[2802] = 2'h3;
    T2[2803] = 2'h0;
    T2[2804] = 2'h2;
    T2[2805] = 2'h1;
    T2[2806] = 2'h0;
    T2[2807] = 2'h3;
    T2[2808] = 2'h0;
    T2[2809] = 2'h2;
    T2[2810] = 2'h2;
    T2[2811] = 2'h0;
    T2[2812] = 2'h3;
    T2[2813] = 2'h0;
    T2[2814] = 2'h2;
    T2[2815] = 2'h3;
    T2[2816] = 2'h0;
    T2[2817] = 2'h3;
    T2[2818] = 2'h0;
    T2[2819] = 2'h2;
    T2[2820] = 2'h0;
    T2[2821] = 2'h1;
    T2[2822] = 2'h3;
    T2[2823] = 2'h0;
    T2[2824] = 2'h2;
    T2[2825] = 2'h1;
    T2[2826] = 2'h1;
    T2[2827] = 2'h3;
    T2[2828] = 2'h0;
    T2[2829] = 2'h2;
    T2[2830] = 2'h2;
    T2[2831] = 2'h1;
    T2[2832] = 2'h3;
    T2[2833] = 2'h0;
    T2[2834] = 2'h2;
    T2[2835] = 2'h3;
    T2[2836] = 2'h1;
    T2[2837] = 2'h3;
    T2[2838] = 2'h0;
    T2[2839] = 2'h2;
    T2[2840] = 2'h0;
    T2[2841] = 2'h2;
    T2[2842] = 2'h3;
    T2[2843] = 2'h0;
    T2[2844] = 2'h2;
    T2[2845] = 2'h1;
    T2[2846] = 2'h2;
    T2[2847] = 2'h3;
    T2[2848] = 2'h0;
    T2[2849] = 2'h2;
    T2[2850] = 2'h2;
    T2[2851] = 2'h2;
    T2[2852] = 2'h3;
    T2[2853] = 2'h0;
    T2[2854] = 2'h2;
    T2[2855] = 2'h3;
    T2[2856] = 2'h2;
    T2[2857] = 2'h3;
    T2[2858] = 2'h0;
    T2[2859] = 2'h2;
    T2[2860] = 2'h0;
    T2[2861] = 2'h3;
    T2[2862] = 2'h3;
    T2[2863] = 2'h0;
    T2[2864] = 2'h2;
    T2[2865] = 2'h1;
    T2[2866] = 2'h3;
    T2[2867] = 2'h3;
    T2[2868] = 2'h0;
    T2[2869] = 2'h2;
    T2[2870] = 2'h2;
    T2[2871] = 2'h3;
    T2[2872] = 2'h3;
    T2[2873] = 2'h0;
    T2[2874] = 2'h2;
    T2[2875] = 2'h3;
    T2[2876] = 2'h3;
    T2[2877] = 2'h3;
    T2[2878] = 2'h0;
    T2[2879] = 2'h2;
    T2[2880] = 2'h0;
    T2[2881] = 2'h0;
    T2[2882] = 2'h0;
    T2[2883] = 2'h1;
    T2[2884] = 2'h2;
    T2[2885] = 2'h1;
    T2[2886] = 2'h0;
    T2[2887] = 2'h0;
    T2[2888] = 2'h1;
    T2[2889] = 2'h2;
    T2[2890] = 2'h2;
    T2[2891] = 2'h0;
    T2[2892] = 2'h0;
    T2[2893] = 2'h1;
    T2[2894] = 2'h2;
    T2[2895] = 2'h3;
    T2[2896] = 2'h0;
    T2[2897] = 2'h0;
    T2[2898] = 2'h1;
    T2[2899] = 2'h2;
    T2[2900] = 2'h0;
    T2[2901] = 2'h1;
    T2[2902] = 2'h0;
    T2[2903] = 2'h1;
    T2[2904] = 2'h2;
    T2[2905] = 2'h1;
    T2[2906] = 2'h1;
    T2[2907] = 2'h0;
    T2[2908] = 2'h1;
    T2[2909] = 2'h2;
    T2[2910] = 2'h2;
    T2[2911] = 2'h1;
    T2[2912] = 2'h0;
    T2[2913] = 2'h1;
    T2[2914] = 2'h2;
    T2[2915] = 2'h3;
    T2[2916] = 2'h1;
    T2[2917] = 2'h0;
    T2[2918] = 2'h1;
    T2[2919] = 2'h2;
    T2[2920] = 2'h0;
    T2[2921] = 2'h2;
    T2[2922] = 2'h0;
    T2[2923] = 2'h1;
    T2[2924] = 2'h2;
    T2[2925] = 2'h1;
    T2[2926] = 2'h2;
    T2[2927] = 2'h0;
    T2[2928] = 2'h1;
    T2[2929] = 2'h2;
    T2[2930] = 2'h2;
    T2[2931] = 2'h2;
    T2[2932] = 2'h0;
    T2[2933] = 2'h1;
    T2[2934] = 2'h2;
    T2[2935] = 2'h3;
    T2[2936] = 2'h2;
    T2[2937] = 2'h0;
    T2[2938] = 2'h1;
    T2[2939] = 2'h2;
    T2[2940] = 2'h0;
    T2[2941] = 2'h3;
    T2[2942] = 2'h0;
    T2[2943] = 2'h1;
    T2[2944] = 2'h2;
    T2[2945] = 2'h1;
    T2[2946] = 2'h3;
    T2[2947] = 2'h0;
    T2[2948] = 2'h1;
    T2[2949] = 2'h2;
    T2[2950] = 2'h2;
    T2[2951] = 2'h3;
    T2[2952] = 2'h0;
    T2[2953] = 2'h1;
    T2[2954] = 2'h2;
    T2[2955] = 2'h3;
    T2[2956] = 2'h3;
    T2[2957] = 2'h0;
    T2[2958] = 2'h1;
    T2[2959] = 2'h2;
    T2[2960] = 2'h0;
    T2[2961] = 2'h0;
    T2[2962] = 2'h1;
    T2[2963] = 2'h1;
    T2[2964] = 2'h2;
    T2[2965] = 2'h1;
    T2[2966] = 2'h0;
    T2[2967] = 2'h1;
    T2[2968] = 2'h1;
    T2[2969] = 2'h2;
    T2[2970] = 2'h2;
    T2[2971] = 2'h0;
    T2[2972] = 2'h1;
    T2[2973] = 2'h1;
    T2[2974] = 2'h2;
    T2[2975] = 2'h3;
    T2[2976] = 2'h0;
    T2[2977] = 2'h1;
    T2[2978] = 2'h1;
    T2[2979] = 2'h2;
    T2[2980] = 2'h0;
    T2[2981] = 2'h1;
    T2[2982] = 2'h1;
    T2[2983] = 2'h1;
    T2[2984] = 2'h2;
    T2[2985] = 2'h1;
    T2[2986] = 2'h1;
    T2[2987] = 2'h1;
    T2[2988] = 2'h1;
    T2[2989] = 2'h2;
    T2[2990] = 2'h2;
    T2[2991] = 2'h1;
    T2[2992] = 2'h1;
    T2[2993] = 2'h1;
    T2[2994] = 2'h2;
    T2[2995] = 2'h3;
    T2[2996] = 2'h1;
    T2[2997] = 2'h1;
    T2[2998] = 2'h1;
    T2[2999] = 2'h2;
    T2[3000] = 2'h0;
    T2[3001] = 2'h2;
    T2[3002] = 2'h1;
    T2[3003] = 2'h1;
    T2[3004] = 2'h2;
    T2[3005] = 2'h1;
    T2[3006] = 2'h2;
    T2[3007] = 2'h1;
    T2[3008] = 2'h1;
    T2[3009] = 2'h2;
    T2[3010] = 2'h2;
    T2[3011] = 2'h2;
    T2[3012] = 2'h1;
    T2[3013] = 2'h1;
    T2[3014] = 2'h2;
    T2[3015] = 2'h3;
    T2[3016] = 2'h2;
    T2[3017] = 2'h1;
    T2[3018] = 2'h1;
    T2[3019] = 2'h2;
    T2[3020] = 2'h0;
    T2[3021] = 2'h3;
    T2[3022] = 2'h1;
    T2[3023] = 2'h1;
    T2[3024] = 2'h2;
    T2[3025] = 2'h1;
    T2[3026] = 2'h3;
    T2[3027] = 2'h1;
    T2[3028] = 2'h1;
    T2[3029] = 2'h2;
    T2[3030] = 2'h2;
    T2[3031] = 2'h3;
    T2[3032] = 2'h1;
    T2[3033] = 2'h1;
    T2[3034] = 2'h2;
    T2[3035] = 2'h3;
    T2[3036] = 2'h3;
    T2[3037] = 2'h1;
    T2[3038] = 2'h1;
    T2[3039] = 2'h2;
    T2[3040] = 2'h0;
    T2[3041] = 2'h0;
    T2[3042] = 2'h2;
    T2[3043] = 2'h1;
    T2[3044] = 2'h2;
    T2[3045] = 2'h1;
    T2[3046] = 2'h0;
    T2[3047] = 2'h2;
    T2[3048] = 2'h1;
    T2[3049] = 2'h2;
    T2[3050] = 2'h2;
    T2[3051] = 2'h0;
    T2[3052] = 2'h2;
    T2[3053] = 2'h1;
    T2[3054] = 2'h2;
    T2[3055] = 2'h3;
    T2[3056] = 2'h0;
    T2[3057] = 2'h2;
    T2[3058] = 2'h1;
    T2[3059] = 2'h2;
    T2[3060] = 2'h0;
    T2[3061] = 2'h1;
    T2[3062] = 2'h2;
    T2[3063] = 2'h1;
    T2[3064] = 2'h2;
    T2[3065] = 2'h1;
    T2[3066] = 2'h1;
    T2[3067] = 2'h2;
    T2[3068] = 2'h1;
    T2[3069] = 2'h2;
    T2[3070] = 2'h2;
    T2[3071] = 2'h1;
    T2[3072] = 2'h2;
    T2[3073] = 2'h1;
    T2[3074] = 2'h2;
    T2[3075] = 2'h3;
    T2[3076] = 2'h1;
    T2[3077] = 2'h2;
    T2[3078] = 2'h1;
    T2[3079] = 2'h2;
    T2[3080] = 2'h0;
    T2[3081] = 2'h2;
    T2[3082] = 2'h2;
    T2[3083] = 2'h1;
    T2[3084] = 2'h2;
    T2[3085] = 2'h1;
    T2[3086] = 2'h2;
    T2[3087] = 2'h2;
    T2[3088] = 2'h1;
    T2[3089] = 2'h2;
    T2[3090] = 2'h2;
    T2[3091] = 2'h2;
    T2[3092] = 2'h2;
    T2[3093] = 2'h1;
    T2[3094] = 2'h2;
    T2[3095] = 2'h3;
    T2[3096] = 2'h2;
    T2[3097] = 2'h2;
    T2[3098] = 2'h1;
    T2[3099] = 2'h2;
    T2[3100] = 2'h0;
    T2[3101] = 2'h3;
    T2[3102] = 2'h2;
    T2[3103] = 2'h1;
    T2[3104] = 2'h2;
    T2[3105] = 2'h1;
    T2[3106] = 2'h3;
    T2[3107] = 2'h2;
    T2[3108] = 2'h1;
    T2[3109] = 2'h2;
    T2[3110] = 2'h2;
    T2[3111] = 2'h3;
    T2[3112] = 2'h2;
    T2[3113] = 2'h1;
    T2[3114] = 2'h2;
    T2[3115] = 2'h3;
    T2[3116] = 2'h3;
    T2[3117] = 2'h2;
    T2[3118] = 2'h1;
    T2[3119] = 2'h2;
    T2[3120] = 2'h0;
    T2[3121] = 2'h0;
    T2[3122] = 2'h3;
    T2[3123] = 2'h1;
    T2[3124] = 2'h2;
    T2[3125] = 2'h1;
    T2[3126] = 2'h0;
    T2[3127] = 2'h3;
    T2[3128] = 2'h1;
    T2[3129] = 2'h2;
    T2[3130] = 2'h2;
    T2[3131] = 2'h0;
    T2[3132] = 2'h3;
    T2[3133] = 2'h1;
    T2[3134] = 2'h2;
    T2[3135] = 2'h3;
    T2[3136] = 2'h0;
    T2[3137] = 2'h3;
    T2[3138] = 2'h1;
    T2[3139] = 2'h2;
    T2[3140] = 2'h0;
    T2[3141] = 2'h1;
    T2[3142] = 2'h3;
    T2[3143] = 2'h1;
    T2[3144] = 2'h2;
    T2[3145] = 2'h1;
    T2[3146] = 2'h1;
    T2[3147] = 2'h3;
    T2[3148] = 2'h1;
    T2[3149] = 2'h2;
    T2[3150] = 2'h2;
    T2[3151] = 2'h1;
    T2[3152] = 2'h3;
    T2[3153] = 2'h1;
    T2[3154] = 2'h2;
    T2[3155] = 2'h3;
    T2[3156] = 2'h1;
    T2[3157] = 2'h3;
    T2[3158] = 2'h1;
    T2[3159] = 2'h2;
    T2[3160] = 2'h0;
    T2[3161] = 2'h2;
    T2[3162] = 2'h3;
    T2[3163] = 2'h1;
    T2[3164] = 2'h2;
    T2[3165] = 2'h1;
    T2[3166] = 2'h2;
    T2[3167] = 2'h3;
    T2[3168] = 2'h1;
    T2[3169] = 2'h2;
    T2[3170] = 2'h2;
    T2[3171] = 2'h2;
    T2[3172] = 2'h3;
    T2[3173] = 2'h1;
    T2[3174] = 2'h2;
    T2[3175] = 2'h3;
    T2[3176] = 2'h2;
    T2[3177] = 2'h3;
    T2[3178] = 2'h1;
    T2[3179] = 2'h2;
    T2[3180] = 2'h0;
    T2[3181] = 2'h3;
    T2[3182] = 2'h3;
    T2[3183] = 2'h1;
    T2[3184] = 2'h2;
    T2[3185] = 2'h1;
    T2[3186] = 2'h3;
    T2[3187] = 2'h3;
    T2[3188] = 2'h1;
    T2[3189] = 2'h2;
    T2[3190] = 2'h2;
    T2[3191] = 2'h3;
    T2[3192] = 2'h3;
    T2[3193] = 2'h1;
    T2[3194] = 2'h2;
    T2[3195] = 2'h3;
    T2[3196] = 2'h3;
    T2[3197] = 2'h3;
    T2[3198] = 2'h1;
    T2[3199] = 2'h2;
    T2[3200] = 2'h0;
    T2[3201] = 2'h0;
    T2[3202] = 2'h0;
    T2[3203] = 2'h2;
    T2[3204] = 2'h2;
    T2[3205] = 2'h1;
    T2[3206] = 2'h0;
    T2[3207] = 2'h0;
    T2[3208] = 2'h2;
    T2[3209] = 2'h2;
    T2[3210] = 2'h2;
    T2[3211] = 2'h0;
    T2[3212] = 2'h0;
    T2[3213] = 2'h2;
    T2[3214] = 2'h2;
    T2[3215] = 2'h3;
    T2[3216] = 2'h0;
    T2[3217] = 2'h0;
    T2[3218] = 2'h2;
    T2[3219] = 2'h2;
    T2[3220] = 2'h0;
    T2[3221] = 2'h1;
    T2[3222] = 2'h0;
    T2[3223] = 2'h2;
    T2[3224] = 2'h2;
    T2[3225] = 2'h1;
    T2[3226] = 2'h1;
    T2[3227] = 2'h0;
    T2[3228] = 2'h2;
    T2[3229] = 2'h2;
    T2[3230] = 2'h2;
    T2[3231] = 2'h1;
    T2[3232] = 2'h0;
    T2[3233] = 2'h2;
    T2[3234] = 2'h2;
    T2[3235] = 2'h3;
    T2[3236] = 2'h1;
    T2[3237] = 2'h0;
    T2[3238] = 2'h2;
    T2[3239] = 2'h2;
    T2[3240] = 2'h0;
    T2[3241] = 2'h2;
    T2[3242] = 2'h0;
    T2[3243] = 2'h2;
    T2[3244] = 2'h2;
    T2[3245] = 2'h1;
    T2[3246] = 2'h2;
    T2[3247] = 2'h0;
    T2[3248] = 2'h2;
    T2[3249] = 2'h2;
    T2[3250] = 2'h2;
    T2[3251] = 2'h2;
    T2[3252] = 2'h0;
    T2[3253] = 2'h2;
    T2[3254] = 2'h2;
    T2[3255] = 2'h3;
    T2[3256] = 2'h2;
    T2[3257] = 2'h0;
    T2[3258] = 2'h2;
    T2[3259] = 2'h2;
    T2[3260] = 2'h0;
    T2[3261] = 2'h3;
    T2[3262] = 2'h0;
    T2[3263] = 2'h2;
    T2[3264] = 2'h2;
    T2[3265] = 2'h1;
    T2[3266] = 2'h3;
    T2[3267] = 2'h0;
    T2[3268] = 2'h2;
    T2[3269] = 2'h2;
    T2[3270] = 2'h2;
    T2[3271] = 2'h3;
    T2[3272] = 2'h0;
    T2[3273] = 2'h2;
    T2[3274] = 2'h2;
    T2[3275] = 2'h3;
    T2[3276] = 2'h3;
    T2[3277] = 2'h0;
    T2[3278] = 2'h2;
    T2[3279] = 2'h2;
    T2[3280] = 2'h0;
    T2[3281] = 2'h0;
    T2[3282] = 2'h1;
    T2[3283] = 2'h2;
    T2[3284] = 2'h2;
    T2[3285] = 2'h1;
    T2[3286] = 2'h0;
    T2[3287] = 2'h1;
    T2[3288] = 2'h2;
    T2[3289] = 2'h2;
    T2[3290] = 2'h2;
    T2[3291] = 2'h0;
    T2[3292] = 2'h1;
    T2[3293] = 2'h2;
    T2[3294] = 2'h2;
    T2[3295] = 2'h3;
    T2[3296] = 2'h0;
    T2[3297] = 2'h1;
    T2[3298] = 2'h2;
    T2[3299] = 2'h2;
    T2[3300] = 2'h0;
    T2[3301] = 2'h1;
    T2[3302] = 2'h1;
    T2[3303] = 2'h2;
    T2[3304] = 2'h2;
    T2[3305] = 2'h1;
    T2[3306] = 2'h1;
    T2[3307] = 2'h1;
    T2[3308] = 2'h2;
    T2[3309] = 2'h2;
    T2[3310] = 2'h2;
    T2[3311] = 2'h1;
    T2[3312] = 2'h1;
    T2[3313] = 2'h2;
    T2[3314] = 2'h2;
    T2[3315] = 2'h3;
    T2[3316] = 2'h1;
    T2[3317] = 2'h1;
    T2[3318] = 2'h2;
    T2[3319] = 2'h2;
    T2[3320] = 2'h0;
    T2[3321] = 2'h2;
    T2[3322] = 2'h1;
    T2[3323] = 2'h2;
    T2[3324] = 2'h2;
    T2[3325] = 2'h1;
    T2[3326] = 2'h2;
    T2[3327] = 2'h1;
    T2[3328] = 2'h2;
    T2[3329] = 2'h2;
    T2[3330] = 2'h2;
    T2[3331] = 2'h2;
    T2[3332] = 2'h1;
    T2[3333] = 2'h2;
    T2[3334] = 2'h2;
    T2[3335] = 2'h3;
    T2[3336] = 2'h2;
    T2[3337] = 2'h1;
    T2[3338] = 2'h2;
    T2[3339] = 2'h2;
    T2[3340] = 2'h0;
    T2[3341] = 2'h3;
    T2[3342] = 2'h1;
    T2[3343] = 2'h2;
    T2[3344] = 2'h2;
    T2[3345] = 2'h1;
    T2[3346] = 2'h3;
    T2[3347] = 2'h1;
    T2[3348] = 2'h2;
    T2[3349] = 2'h2;
    T2[3350] = 2'h2;
    T2[3351] = 2'h3;
    T2[3352] = 2'h1;
    T2[3353] = 2'h2;
    T2[3354] = 2'h2;
    T2[3355] = 2'h3;
    T2[3356] = 2'h3;
    T2[3357] = 2'h1;
    T2[3358] = 2'h2;
    T2[3359] = 2'h2;
    T2[3360] = 2'h0;
    T2[3361] = 2'h0;
    T2[3362] = 2'h2;
    T2[3363] = 2'h2;
    T2[3364] = 2'h2;
    T2[3365] = 2'h1;
    T2[3366] = 2'h0;
    T2[3367] = 2'h2;
    T2[3368] = 2'h2;
    T2[3369] = 2'h2;
    T2[3370] = 2'h2;
    T2[3371] = 2'h0;
    T2[3372] = 2'h2;
    T2[3373] = 2'h2;
    T2[3374] = 2'h2;
    T2[3375] = 2'h3;
    T2[3376] = 2'h0;
    T2[3377] = 2'h2;
    T2[3378] = 2'h2;
    T2[3379] = 2'h2;
    T2[3380] = 2'h0;
    T2[3381] = 2'h1;
    T2[3382] = 2'h2;
    T2[3383] = 2'h2;
    T2[3384] = 2'h2;
    T2[3385] = 2'h1;
    T2[3386] = 2'h1;
    T2[3387] = 2'h2;
    T2[3388] = 2'h2;
    T2[3389] = 2'h2;
    T2[3390] = 2'h2;
    T2[3391] = 2'h1;
    T2[3392] = 2'h2;
    T2[3393] = 2'h2;
    T2[3394] = 2'h2;
    T2[3395] = 2'h3;
    T2[3396] = 2'h1;
    T2[3397] = 2'h2;
    T2[3398] = 2'h2;
    T2[3399] = 2'h2;
    T2[3400] = 2'h0;
    T2[3401] = 2'h2;
    T2[3402] = 2'h2;
    T2[3403] = 2'h2;
    T2[3404] = 2'h2;
    T2[3405] = 2'h1;
    T2[3406] = 2'h2;
    T2[3407] = 2'h2;
    T2[3408] = 2'h2;
    T2[3409] = 2'h2;
    T2[3410] = 2'h2;
    T2[3411] = 2'h2;
    T2[3412] = 2'h2;
    T2[3413] = 2'h2;
    T2[3414] = 2'h2;
    T2[3415] = 2'h3;
    T2[3416] = 2'h2;
    T2[3417] = 2'h2;
    T2[3418] = 2'h2;
    T2[3419] = 2'h2;
    T2[3420] = 2'h0;
    T2[3421] = 2'h3;
    T2[3422] = 2'h2;
    T2[3423] = 2'h2;
    T2[3424] = 2'h2;
    T2[3425] = 2'h1;
    T2[3426] = 2'h3;
    T2[3427] = 2'h2;
    T2[3428] = 2'h2;
    T2[3429] = 2'h2;
    T2[3430] = 2'h2;
    T2[3431] = 2'h3;
    T2[3432] = 2'h2;
    T2[3433] = 2'h2;
    T2[3434] = 2'h2;
    T2[3435] = 2'h3;
    T2[3436] = 2'h3;
    T2[3437] = 2'h2;
    T2[3438] = 2'h2;
    T2[3439] = 2'h2;
    T2[3440] = 2'h0;
    T2[3441] = 2'h0;
    T2[3442] = 2'h3;
    T2[3443] = 2'h2;
    T2[3444] = 2'h2;
    T2[3445] = 2'h1;
    T2[3446] = 2'h0;
    T2[3447] = 2'h3;
    T2[3448] = 2'h2;
    T2[3449] = 2'h2;
    T2[3450] = 2'h2;
    T2[3451] = 2'h0;
    T2[3452] = 2'h3;
    T2[3453] = 2'h2;
    T2[3454] = 2'h2;
    T2[3455] = 2'h3;
    T2[3456] = 2'h0;
    T2[3457] = 2'h3;
    T2[3458] = 2'h2;
    T2[3459] = 2'h2;
    T2[3460] = 2'h0;
    T2[3461] = 2'h1;
    T2[3462] = 2'h3;
    T2[3463] = 2'h2;
    T2[3464] = 2'h2;
    T2[3465] = 2'h1;
    T2[3466] = 2'h1;
    T2[3467] = 2'h3;
    T2[3468] = 2'h2;
    T2[3469] = 2'h2;
    T2[3470] = 2'h2;
    T2[3471] = 2'h1;
    T2[3472] = 2'h3;
    T2[3473] = 2'h2;
    T2[3474] = 2'h2;
    T2[3475] = 2'h3;
    T2[3476] = 2'h1;
    T2[3477] = 2'h3;
    T2[3478] = 2'h2;
    T2[3479] = 2'h2;
    T2[3480] = 2'h0;
    T2[3481] = 2'h2;
    T2[3482] = 2'h3;
    T2[3483] = 2'h2;
    T2[3484] = 2'h2;
    T2[3485] = 2'h1;
    T2[3486] = 2'h2;
    T2[3487] = 2'h3;
    T2[3488] = 2'h2;
    T2[3489] = 2'h2;
    T2[3490] = 2'h2;
    T2[3491] = 2'h2;
    T2[3492] = 2'h3;
    T2[3493] = 2'h2;
    T2[3494] = 2'h2;
    T2[3495] = 2'h3;
    T2[3496] = 2'h2;
    T2[3497] = 2'h3;
    T2[3498] = 2'h2;
    T2[3499] = 2'h2;
    T2[3500] = 2'h0;
    T2[3501] = 2'h3;
    T2[3502] = 2'h3;
    T2[3503] = 2'h2;
    T2[3504] = 2'h2;
    T2[3505] = 2'h1;
    T2[3506] = 2'h3;
    T2[3507] = 2'h3;
    T2[3508] = 2'h2;
    T2[3509] = 2'h2;
    T2[3510] = 2'h2;
    T2[3511] = 2'h3;
    T2[3512] = 2'h3;
    T2[3513] = 2'h2;
    T2[3514] = 2'h2;
    T2[3515] = 2'h3;
    T2[3516] = 2'h3;
    T2[3517] = 2'h3;
    T2[3518] = 2'h2;
    T2[3519] = 2'h2;
    T2[3520] = 2'h0;
    T2[3521] = 2'h0;
    T2[3522] = 2'h0;
    T2[3523] = 2'h3;
    T2[3524] = 2'h2;
    T2[3525] = 2'h1;
    T2[3526] = 2'h0;
    T2[3527] = 2'h0;
    T2[3528] = 2'h3;
    T2[3529] = 2'h2;
    T2[3530] = 2'h2;
    T2[3531] = 2'h0;
    T2[3532] = 2'h0;
    T2[3533] = 2'h3;
    T2[3534] = 2'h2;
    T2[3535] = 2'h3;
    T2[3536] = 2'h0;
    T2[3537] = 2'h0;
    T2[3538] = 2'h3;
    T2[3539] = 2'h2;
    T2[3540] = 2'h0;
    T2[3541] = 2'h1;
    T2[3542] = 2'h0;
    T2[3543] = 2'h3;
    T2[3544] = 2'h2;
    T2[3545] = 2'h1;
    T2[3546] = 2'h1;
    T2[3547] = 2'h0;
    T2[3548] = 2'h3;
    T2[3549] = 2'h2;
    T2[3550] = 2'h2;
    T2[3551] = 2'h1;
    T2[3552] = 2'h0;
    T2[3553] = 2'h3;
    T2[3554] = 2'h2;
    T2[3555] = 2'h3;
    T2[3556] = 2'h1;
    T2[3557] = 2'h0;
    T2[3558] = 2'h3;
    T2[3559] = 2'h2;
    T2[3560] = 2'h0;
    T2[3561] = 2'h2;
    T2[3562] = 2'h0;
    T2[3563] = 2'h3;
    T2[3564] = 2'h2;
    T2[3565] = 2'h1;
    T2[3566] = 2'h2;
    T2[3567] = 2'h0;
    T2[3568] = 2'h3;
    T2[3569] = 2'h2;
    T2[3570] = 2'h2;
    T2[3571] = 2'h2;
    T2[3572] = 2'h0;
    T2[3573] = 2'h3;
    T2[3574] = 2'h2;
    T2[3575] = 2'h3;
    T2[3576] = 2'h2;
    T2[3577] = 2'h0;
    T2[3578] = 2'h3;
    T2[3579] = 2'h2;
    T2[3580] = 2'h0;
    T2[3581] = 2'h3;
    T2[3582] = 2'h0;
    T2[3583] = 2'h3;
    T2[3584] = 2'h2;
    T2[3585] = 2'h1;
    T2[3586] = 2'h3;
    T2[3587] = 2'h0;
    T2[3588] = 2'h3;
    T2[3589] = 2'h2;
    T2[3590] = 2'h2;
    T2[3591] = 2'h3;
    T2[3592] = 2'h0;
    T2[3593] = 2'h3;
    T2[3594] = 2'h2;
    T2[3595] = 2'h3;
    T2[3596] = 2'h3;
    T2[3597] = 2'h0;
    T2[3598] = 2'h3;
    T2[3599] = 2'h2;
    T2[3600] = 2'h0;
    T2[3601] = 2'h0;
    T2[3602] = 2'h1;
    T2[3603] = 2'h3;
    T2[3604] = 2'h2;
    T2[3605] = 2'h1;
    T2[3606] = 2'h0;
    T2[3607] = 2'h1;
    T2[3608] = 2'h3;
    T2[3609] = 2'h2;
    T2[3610] = 2'h2;
    T2[3611] = 2'h0;
    T2[3612] = 2'h1;
    T2[3613] = 2'h3;
    T2[3614] = 2'h2;
    T2[3615] = 2'h3;
    T2[3616] = 2'h0;
    T2[3617] = 2'h1;
    T2[3618] = 2'h3;
    T2[3619] = 2'h2;
    T2[3620] = 2'h0;
    T2[3621] = 2'h1;
    T2[3622] = 2'h1;
    T2[3623] = 2'h3;
    T2[3624] = 2'h2;
    T2[3625] = 2'h1;
    T2[3626] = 2'h1;
    T2[3627] = 2'h1;
    T2[3628] = 2'h3;
    T2[3629] = 2'h2;
    T2[3630] = 2'h2;
    T2[3631] = 2'h1;
    T2[3632] = 2'h1;
    T2[3633] = 2'h3;
    T2[3634] = 2'h2;
    T2[3635] = 2'h3;
    T2[3636] = 2'h1;
    T2[3637] = 2'h1;
    T2[3638] = 2'h3;
    T2[3639] = 2'h2;
    T2[3640] = 2'h0;
    T2[3641] = 2'h2;
    T2[3642] = 2'h1;
    T2[3643] = 2'h3;
    T2[3644] = 2'h2;
    T2[3645] = 2'h1;
    T2[3646] = 2'h2;
    T2[3647] = 2'h1;
    T2[3648] = 2'h3;
    T2[3649] = 2'h2;
    T2[3650] = 2'h2;
    T2[3651] = 2'h2;
    T2[3652] = 2'h1;
    T2[3653] = 2'h3;
    T2[3654] = 2'h2;
    T2[3655] = 2'h3;
    T2[3656] = 2'h2;
    T2[3657] = 2'h1;
    T2[3658] = 2'h3;
    T2[3659] = 2'h2;
    T2[3660] = 2'h0;
    T2[3661] = 2'h3;
    T2[3662] = 2'h1;
    T2[3663] = 2'h3;
    T2[3664] = 2'h2;
    T2[3665] = 2'h1;
    T2[3666] = 2'h3;
    T2[3667] = 2'h1;
    T2[3668] = 2'h3;
    T2[3669] = 2'h2;
    T2[3670] = 2'h2;
    T2[3671] = 2'h3;
    T2[3672] = 2'h1;
    T2[3673] = 2'h3;
    T2[3674] = 2'h2;
    T2[3675] = 2'h3;
    T2[3676] = 2'h3;
    T2[3677] = 2'h1;
    T2[3678] = 2'h3;
    T2[3679] = 2'h2;
    T2[3680] = 2'h0;
    T2[3681] = 2'h0;
    T2[3682] = 2'h2;
    T2[3683] = 2'h3;
    T2[3684] = 2'h2;
    T2[3685] = 2'h1;
    T2[3686] = 2'h0;
    T2[3687] = 2'h2;
    T2[3688] = 2'h3;
    T2[3689] = 2'h2;
    T2[3690] = 2'h2;
    T2[3691] = 2'h0;
    T2[3692] = 2'h2;
    T2[3693] = 2'h3;
    T2[3694] = 2'h2;
    T2[3695] = 2'h3;
    T2[3696] = 2'h0;
    T2[3697] = 2'h2;
    T2[3698] = 2'h3;
    T2[3699] = 2'h2;
    T2[3700] = 2'h0;
    T2[3701] = 2'h1;
    T2[3702] = 2'h2;
    T2[3703] = 2'h3;
    T2[3704] = 2'h2;
    T2[3705] = 2'h1;
    T2[3706] = 2'h1;
    T2[3707] = 2'h2;
    T2[3708] = 2'h3;
    T2[3709] = 2'h2;
    T2[3710] = 2'h2;
    T2[3711] = 2'h1;
    T2[3712] = 2'h2;
    T2[3713] = 2'h3;
    T2[3714] = 2'h2;
    T2[3715] = 2'h3;
    T2[3716] = 2'h1;
    T2[3717] = 2'h2;
    T2[3718] = 2'h3;
    T2[3719] = 2'h2;
    T2[3720] = 2'h0;
    T2[3721] = 2'h2;
    T2[3722] = 2'h2;
    T2[3723] = 2'h3;
    T2[3724] = 2'h2;
    T2[3725] = 2'h1;
    T2[3726] = 2'h2;
    T2[3727] = 2'h2;
    T2[3728] = 2'h3;
    T2[3729] = 2'h2;
    T2[3730] = 2'h2;
    T2[3731] = 2'h2;
    T2[3732] = 2'h2;
    T2[3733] = 2'h3;
    T2[3734] = 2'h2;
    T2[3735] = 2'h3;
    T2[3736] = 2'h2;
    T2[3737] = 2'h2;
    T2[3738] = 2'h3;
    T2[3739] = 2'h2;
    T2[3740] = 2'h0;
    T2[3741] = 2'h3;
    T2[3742] = 2'h2;
    T2[3743] = 2'h3;
    T2[3744] = 2'h2;
    T2[3745] = 2'h1;
    T2[3746] = 2'h3;
    T2[3747] = 2'h2;
    T2[3748] = 2'h3;
    T2[3749] = 2'h2;
    T2[3750] = 2'h2;
    T2[3751] = 2'h3;
    T2[3752] = 2'h2;
    T2[3753] = 2'h3;
    T2[3754] = 2'h2;
    T2[3755] = 2'h3;
    T2[3756] = 2'h3;
    T2[3757] = 2'h2;
    T2[3758] = 2'h3;
    T2[3759] = 2'h2;
    T2[3760] = 2'h0;
    T2[3761] = 2'h0;
    T2[3762] = 2'h3;
    T2[3763] = 2'h3;
    T2[3764] = 2'h2;
    T2[3765] = 2'h1;
    T2[3766] = 2'h0;
    T2[3767] = 2'h3;
    T2[3768] = 2'h3;
    T2[3769] = 2'h2;
    T2[3770] = 2'h2;
    T2[3771] = 2'h0;
    T2[3772] = 2'h3;
    T2[3773] = 2'h3;
    T2[3774] = 2'h2;
    T2[3775] = 2'h3;
    T2[3776] = 2'h0;
    T2[3777] = 2'h3;
    T2[3778] = 2'h3;
    T2[3779] = 2'h2;
    T2[3780] = 2'h0;
    T2[3781] = 2'h1;
    T2[3782] = 2'h3;
    T2[3783] = 2'h3;
    T2[3784] = 2'h2;
    T2[3785] = 2'h1;
    T2[3786] = 2'h1;
    T2[3787] = 2'h3;
    T2[3788] = 2'h3;
    T2[3789] = 2'h2;
    T2[3790] = 2'h2;
    T2[3791] = 2'h1;
    T2[3792] = 2'h3;
    T2[3793] = 2'h3;
    T2[3794] = 2'h2;
    T2[3795] = 2'h3;
    T2[3796] = 2'h1;
    T2[3797] = 2'h3;
    T2[3798] = 2'h3;
    T2[3799] = 2'h2;
    T2[3800] = 2'h0;
    T2[3801] = 2'h2;
    T2[3802] = 2'h3;
    T2[3803] = 2'h3;
    T2[3804] = 2'h2;
    T2[3805] = 2'h1;
    T2[3806] = 2'h2;
    T2[3807] = 2'h3;
    T2[3808] = 2'h3;
    T2[3809] = 2'h2;
    T2[3810] = 2'h2;
    T2[3811] = 2'h2;
    T2[3812] = 2'h3;
    T2[3813] = 2'h3;
    T2[3814] = 2'h2;
    T2[3815] = 2'h3;
    T2[3816] = 2'h2;
    T2[3817] = 2'h3;
    T2[3818] = 2'h3;
    T2[3819] = 2'h2;
    T2[3820] = 2'h0;
    T2[3821] = 2'h3;
    T2[3822] = 2'h3;
    T2[3823] = 2'h3;
    T2[3824] = 2'h2;
    T2[3825] = 2'h1;
    T2[3826] = 2'h3;
    T2[3827] = 2'h3;
    T2[3828] = 2'h3;
    T2[3829] = 2'h2;
    T2[3830] = 2'h2;
    T2[3831] = 2'h3;
    T2[3832] = 2'h3;
    T2[3833] = 2'h3;
    T2[3834] = 2'h2;
    T2[3835] = 2'h3;
    T2[3836] = 2'h3;
    T2[3837] = 2'h3;
    T2[3838] = 2'h3;
    T2[3839] = 2'h2;
    T2[3840] = 2'h0;
    T2[3841] = 2'h0;
    T2[3842] = 2'h0;
    T2[3843] = 2'h0;
    T2[3844] = 2'h3;
    T2[3845] = 2'h1;
    T2[3846] = 2'h0;
    T2[3847] = 2'h0;
    T2[3848] = 2'h0;
    T2[3849] = 2'h3;
    T2[3850] = 2'h2;
    T2[3851] = 2'h0;
    T2[3852] = 2'h0;
    T2[3853] = 2'h0;
    T2[3854] = 2'h3;
    T2[3855] = 2'h3;
    T2[3856] = 2'h0;
    T2[3857] = 2'h0;
    T2[3858] = 2'h0;
    T2[3859] = 2'h3;
    T2[3860] = 2'h0;
    T2[3861] = 2'h1;
    T2[3862] = 2'h0;
    T2[3863] = 2'h0;
    T2[3864] = 2'h3;
    T2[3865] = 2'h1;
    T2[3866] = 2'h1;
    T2[3867] = 2'h0;
    T2[3868] = 2'h0;
    T2[3869] = 2'h3;
    T2[3870] = 2'h2;
    T2[3871] = 2'h1;
    T2[3872] = 2'h0;
    T2[3873] = 2'h0;
    T2[3874] = 2'h3;
    T2[3875] = 2'h3;
    T2[3876] = 2'h1;
    T2[3877] = 2'h0;
    T2[3878] = 2'h0;
    T2[3879] = 2'h3;
    T2[3880] = 2'h0;
    T2[3881] = 2'h2;
    T2[3882] = 2'h0;
    T2[3883] = 2'h0;
    T2[3884] = 2'h3;
    T2[3885] = 2'h1;
    T2[3886] = 2'h2;
    T2[3887] = 2'h0;
    T2[3888] = 2'h0;
    T2[3889] = 2'h3;
    T2[3890] = 2'h2;
    T2[3891] = 2'h2;
    T2[3892] = 2'h0;
    T2[3893] = 2'h0;
    T2[3894] = 2'h3;
    T2[3895] = 2'h3;
    T2[3896] = 2'h2;
    T2[3897] = 2'h0;
    T2[3898] = 2'h0;
    T2[3899] = 2'h3;
    T2[3900] = 2'h0;
    T2[3901] = 2'h3;
    T2[3902] = 2'h0;
    T2[3903] = 2'h0;
    T2[3904] = 2'h3;
    T2[3905] = 2'h1;
    T2[3906] = 2'h3;
    T2[3907] = 2'h0;
    T2[3908] = 2'h0;
    T2[3909] = 2'h3;
    T2[3910] = 2'h2;
    T2[3911] = 2'h3;
    T2[3912] = 2'h0;
    T2[3913] = 2'h0;
    T2[3914] = 2'h3;
    T2[3915] = 2'h3;
    T2[3916] = 2'h3;
    T2[3917] = 2'h0;
    T2[3918] = 2'h0;
    T2[3919] = 2'h3;
    T2[3920] = 2'h0;
    T2[3921] = 2'h0;
    T2[3922] = 2'h1;
    T2[3923] = 2'h0;
    T2[3924] = 2'h3;
    T2[3925] = 2'h1;
    T2[3926] = 2'h0;
    T2[3927] = 2'h1;
    T2[3928] = 2'h0;
    T2[3929] = 2'h3;
    T2[3930] = 2'h2;
    T2[3931] = 2'h0;
    T2[3932] = 2'h1;
    T2[3933] = 2'h0;
    T2[3934] = 2'h3;
    T2[3935] = 2'h3;
    T2[3936] = 2'h0;
    T2[3937] = 2'h1;
    T2[3938] = 2'h0;
    T2[3939] = 2'h3;
    T2[3940] = 2'h0;
    T2[3941] = 2'h1;
    T2[3942] = 2'h1;
    T2[3943] = 2'h0;
    T2[3944] = 2'h3;
    T2[3945] = 2'h1;
    T2[3946] = 2'h1;
    T2[3947] = 2'h1;
    T2[3948] = 2'h0;
    T2[3949] = 2'h3;
    T2[3950] = 2'h2;
    T2[3951] = 2'h1;
    T2[3952] = 2'h1;
    T2[3953] = 2'h0;
    T2[3954] = 2'h3;
    T2[3955] = 2'h3;
    T2[3956] = 2'h1;
    T2[3957] = 2'h1;
    T2[3958] = 2'h0;
    T2[3959] = 2'h3;
    T2[3960] = 2'h0;
    T2[3961] = 2'h2;
    T2[3962] = 2'h1;
    T2[3963] = 2'h0;
    T2[3964] = 2'h3;
    T2[3965] = 2'h1;
    T2[3966] = 2'h2;
    T2[3967] = 2'h1;
    T2[3968] = 2'h0;
    T2[3969] = 2'h3;
    T2[3970] = 2'h2;
    T2[3971] = 2'h2;
    T2[3972] = 2'h1;
    T2[3973] = 2'h0;
    T2[3974] = 2'h3;
    T2[3975] = 2'h3;
    T2[3976] = 2'h2;
    T2[3977] = 2'h1;
    T2[3978] = 2'h0;
    T2[3979] = 2'h3;
    T2[3980] = 2'h0;
    T2[3981] = 2'h3;
    T2[3982] = 2'h1;
    T2[3983] = 2'h0;
    T2[3984] = 2'h3;
    T2[3985] = 2'h1;
    T2[3986] = 2'h3;
    T2[3987] = 2'h1;
    T2[3988] = 2'h0;
    T2[3989] = 2'h3;
    T2[3990] = 2'h2;
    T2[3991] = 2'h3;
    T2[3992] = 2'h1;
    T2[3993] = 2'h0;
    T2[3994] = 2'h3;
    T2[3995] = 2'h3;
    T2[3996] = 2'h3;
    T2[3997] = 2'h1;
    T2[3998] = 2'h0;
    T2[3999] = 2'h3;
    T2[4000] = 2'h0;
    T2[4001] = 2'h0;
    T2[4002] = 2'h2;
    T2[4003] = 2'h0;
    T2[4004] = 2'h3;
    T2[4005] = 2'h1;
    T2[4006] = 2'h0;
    T2[4007] = 2'h2;
    T2[4008] = 2'h0;
    T2[4009] = 2'h3;
    T2[4010] = 2'h2;
    T2[4011] = 2'h0;
    T2[4012] = 2'h2;
    T2[4013] = 2'h0;
    T2[4014] = 2'h3;
    T2[4015] = 2'h3;
    T2[4016] = 2'h0;
    T2[4017] = 2'h2;
    T2[4018] = 2'h0;
    T2[4019] = 2'h3;
    T2[4020] = 2'h0;
    T2[4021] = 2'h1;
    T2[4022] = 2'h2;
    T2[4023] = 2'h0;
    T2[4024] = 2'h3;
    T2[4025] = 2'h1;
    T2[4026] = 2'h1;
    T2[4027] = 2'h2;
    T2[4028] = 2'h0;
    T2[4029] = 2'h3;
    T2[4030] = 2'h2;
    T2[4031] = 2'h1;
    T2[4032] = 2'h2;
    T2[4033] = 2'h0;
    T2[4034] = 2'h3;
    T2[4035] = 2'h3;
    T2[4036] = 2'h1;
    T2[4037] = 2'h2;
    T2[4038] = 2'h0;
    T2[4039] = 2'h3;
    T2[4040] = 2'h0;
    T2[4041] = 2'h2;
    T2[4042] = 2'h2;
    T2[4043] = 2'h0;
    T2[4044] = 2'h3;
    T2[4045] = 2'h1;
    T2[4046] = 2'h2;
    T2[4047] = 2'h2;
    T2[4048] = 2'h0;
    T2[4049] = 2'h3;
    T2[4050] = 2'h2;
    T2[4051] = 2'h2;
    T2[4052] = 2'h2;
    T2[4053] = 2'h0;
    T2[4054] = 2'h3;
    T2[4055] = 2'h3;
    T2[4056] = 2'h2;
    T2[4057] = 2'h2;
    T2[4058] = 2'h0;
    T2[4059] = 2'h3;
    T2[4060] = 2'h0;
    T2[4061] = 2'h3;
    T2[4062] = 2'h2;
    T2[4063] = 2'h0;
    T2[4064] = 2'h3;
    T2[4065] = 2'h1;
    T2[4066] = 2'h3;
    T2[4067] = 2'h2;
    T2[4068] = 2'h0;
    T2[4069] = 2'h3;
    T2[4070] = 2'h2;
    T2[4071] = 2'h3;
    T2[4072] = 2'h2;
    T2[4073] = 2'h0;
    T2[4074] = 2'h3;
    T2[4075] = 2'h3;
    T2[4076] = 2'h3;
    T2[4077] = 2'h2;
    T2[4078] = 2'h0;
    T2[4079] = 2'h3;
    T2[4080] = 2'h0;
    T2[4081] = 2'h0;
    T2[4082] = 2'h3;
    T2[4083] = 2'h0;
    T2[4084] = 2'h3;
    T2[4085] = 2'h1;
    T2[4086] = 2'h0;
    T2[4087] = 2'h3;
    T2[4088] = 2'h0;
    T2[4089] = 2'h3;
    T2[4090] = 2'h2;
    T2[4091] = 2'h0;
    T2[4092] = 2'h3;
    T2[4093] = 2'h0;
    T2[4094] = 2'h3;
    T2[4095] = 2'h3;
    T2[4096] = 2'h0;
    T2[4097] = 2'h3;
    T2[4098] = 2'h0;
    T2[4099] = 2'h3;
    T2[4100] = 2'h0;
    T2[4101] = 2'h1;
    T2[4102] = 2'h3;
    T2[4103] = 2'h0;
    T2[4104] = 2'h3;
    T2[4105] = 2'h1;
    T2[4106] = 2'h1;
    T2[4107] = 2'h3;
    T2[4108] = 2'h0;
    T2[4109] = 2'h3;
    T2[4110] = 2'h2;
    T2[4111] = 2'h1;
    T2[4112] = 2'h3;
    T2[4113] = 2'h0;
    T2[4114] = 2'h3;
    T2[4115] = 2'h3;
    T2[4116] = 2'h1;
    T2[4117] = 2'h3;
    T2[4118] = 2'h0;
    T2[4119] = 2'h3;
    T2[4120] = 2'h0;
    T2[4121] = 2'h2;
    T2[4122] = 2'h3;
    T2[4123] = 2'h0;
    T2[4124] = 2'h3;
    T2[4125] = 2'h1;
    T2[4126] = 2'h2;
    T2[4127] = 2'h3;
    T2[4128] = 2'h0;
    T2[4129] = 2'h3;
    T2[4130] = 2'h2;
    T2[4131] = 2'h2;
    T2[4132] = 2'h3;
    T2[4133] = 2'h0;
    T2[4134] = 2'h3;
    T2[4135] = 2'h3;
    T2[4136] = 2'h2;
    T2[4137] = 2'h3;
    T2[4138] = 2'h0;
    T2[4139] = 2'h3;
    T2[4140] = 2'h0;
    T2[4141] = 2'h3;
    T2[4142] = 2'h3;
    T2[4143] = 2'h0;
    T2[4144] = 2'h3;
    T2[4145] = 2'h1;
    T2[4146] = 2'h3;
    T2[4147] = 2'h3;
    T2[4148] = 2'h0;
    T2[4149] = 2'h3;
    T2[4150] = 2'h2;
    T2[4151] = 2'h3;
    T2[4152] = 2'h3;
    T2[4153] = 2'h0;
    T2[4154] = 2'h3;
    T2[4155] = 2'h3;
    T2[4156] = 2'h3;
    T2[4157] = 2'h3;
    T2[4158] = 2'h0;
    T2[4159] = 2'h3;
    T2[4160] = 2'h0;
    T2[4161] = 2'h0;
    T2[4162] = 2'h0;
    T2[4163] = 2'h1;
    T2[4164] = 2'h3;
    T2[4165] = 2'h1;
    T2[4166] = 2'h0;
    T2[4167] = 2'h0;
    T2[4168] = 2'h1;
    T2[4169] = 2'h3;
    T2[4170] = 2'h2;
    T2[4171] = 2'h0;
    T2[4172] = 2'h0;
    T2[4173] = 2'h1;
    T2[4174] = 2'h3;
    T2[4175] = 2'h3;
    T2[4176] = 2'h0;
    T2[4177] = 2'h0;
    T2[4178] = 2'h1;
    T2[4179] = 2'h3;
    T2[4180] = 2'h0;
    T2[4181] = 2'h1;
    T2[4182] = 2'h0;
    T2[4183] = 2'h1;
    T2[4184] = 2'h3;
    T2[4185] = 2'h1;
    T2[4186] = 2'h1;
    T2[4187] = 2'h0;
    T2[4188] = 2'h1;
    T2[4189] = 2'h3;
    T2[4190] = 2'h2;
    T2[4191] = 2'h1;
    T2[4192] = 2'h0;
    T2[4193] = 2'h1;
    T2[4194] = 2'h3;
    T2[4195] = 2'h3;
    T2[4196] = 2'h1;
    T2[4197] = 2'h0;
    T2[4198] = 2'h1;
    T2[4199] = 2'h3;
    T2[4200] = 2'h0;
    T2[4201] = 2'h2;
    T2[4202] = 2'h0;
    T2[4203] = 2'h1;
    T2[4204] = 2'h3;
    T2[4205] = 2'h1;
    T2[4206] = 2'h2;
    T2[4207] = 2'h0;
    T2[4208] = 2'h1;
    T2[4209] = 2'h3;
    T2[4210] = 2'h2;
    T2[4211] = 2'h2;
    T2[4212] = 2'h0;
    T2[4213] = 2'h1;
    T2[4214] = 2'h3;
    T2[4215] = 2'h3;
    T2[4216] = 2'h2;
    T2[4217] = 2'h0;
    T2[4218] = 2'h1;
    T2[4219] = 2'h3;
    T2[4220] = 2'h0;
    T2[4221] = 2'h3;
    T2[4222] = 2'h0;
    T2[4223] = 2'h1;
    T2[4224] = 2'h3;
    T2[4225] = 2'h1;
    T2[4226] = 2'h3;
    T2[4227] = 2'h0;
    T2[4228] = 2'h1;
    T2[4229] = 2'h3;
    T2[4230] = 2'h2;
    T2[4231] = 2'h3;
    T2[4232] = 2'h0;
    T2[4233] = 2'h1;
    T2[4234] = 2'h3;
    T2[4235] = 2'h3;
    T2[4236] = 2'h3;
    T2[4237] = 2'h0;
    T2[4238] = 2'h1;
    T2[4239] = 2'h3;
    T2[4240] = 2'h0;
    T2[4241] = 2'h0;
    T2[4242] = 2'h1;
    T2[4243] = 2'h1;
    T2[4244] = 2'h3;
    T2[4245] = 2'h1;
    T2[4246] = 2'h0;
    T2[4247] = 2'h1;
    T2[4248] = 2'h1;
    T2[4249] = 2'h3;
    T2[4250] = 2'h2;
    T2[4251] = 2'h0;
    T2[4252] = 2'h1;
    T2[4253] = 2'h1;
    T2[4254] = 2'h3;
    T2[4255] = 2'h3;
    T2[4256] = 2'h0;
    T2[4257] = 2'h1;
    T2[4258] = 2'h1;
    T2[4259] = 2'h3;
    T2[4260] = 2'h0;
    T2[4261] = 2'h1;
    T2[4262] = 2'h1;
    T2[4263] = 2'h1;
    T2[4264] = 2'h3;
    T2[4265] = 2'h1;
    T2[4266] = 2'h1;
    T2[4267] = 2'h1;
    T2[4268] = 2'h1;
    T2[4269] = 2'h3;
    T2[4270] = 2'h2;
    T2[4271] = 2'h1;
    T2[4272] = 2'h1;
    T2[4273] = 2'h1;
    T2[4274] = 2'h3;
    T2[4275] = 2'h3;
    T2[4276] = 2'h1;
    T2[4277] = 2'h1;
    T2[4278] = 2'h1;
    T2[4279] = 2'h3;
    T2[4280] = 2'h0;
    T2[4281] = 2'h2;
    T2[4282] = 2'h1;
    T2[4283] = 2'h1;
    T2[4284] = 2'h3;
    T2[4285] = 2'h1;
    T2[4286] = 2'h2;
    T2[4287] = 2'h1;
    T2[4288] = 2'h1;
    T2[4289] = 2'h3;
    T2[4290] = 2'h2;
    T2[4291] = 2'h2;
    T2[4292] = 2'h1;
    T2[4293] = 2'h1;
    T2[4294] = 2'h3;
    T2[4295] = 2'h3;
    T2[4296] = 2'h2;
    T2[4297] = 2'h1;
    T2[4298] = 2'h1;
    T2[4299] = 2'h3;
    T2[4300] = 2'h0;
    T2[4301] = 2'h3;
    T2[4302] = 2'h1;
    T2[4303] = 2'h1;
    T2[4304] = 2'h3;
    T2[4305] = 2'h1;
    T2[4306] = 2'h3;
    T2[4307] = 2'h1;
    T2[4308] = 2'h1;
    T2[4309] = 2'h3;
    T2[4310] = 2'h2;
    T2[4311] = 2'h3;
    T2[4312] = 2'h1;
    T2[4313] = 2'h1;
    T2[4314] = 2'h3;
    T2[4315] = 2'h3;
    T2[4316] = 2'h3;
    T2[4317] = 2'h1;
    T2[4318] = 2'h1;
    T2[4319] = 2'h3;
    T2[4320] = 2'h0;
    T2[4321] = 2'h0;
    T2[4322] = 2'h2;
    T2[4323] = 2'h1;
    T2[4324] = 2'h3;
    T2[4325] = 2'h1;
    T2[4326] = 2'h0;
    T2[4327] = 2'h2;
    T2[4328] = 2'h1;
    T2[4329] = 2'h3;
    T2[4330] = 2'h2;
    T2[4331] = 2'h0;
    T2[4332] = 2'h2;
    T2[4333] = 2'h1;
    T2[4334] = 2'h3;
    T2[4335] = 2'h3;
    T2[4336] = 2'h0;
    T2[4337] = 2'h2;
    T2[4338] = 2'h1;
    T2[4339] = 2'h3;
    T2[4340] = 2'h0;
    T2[4341] = 2'h1;
    T2[4342] = 2'h2;
    T2[4343] = 2'h1;
    T2[4344] = 2'h3;
    T2[4345] = 2'h1;
    T2[4346] = 2'h1;
    T2[4347] = 2'h2;
    T2[4348] = 2'h1;
    T2[4349] = 2'h3;
    T2[4350] = 2'h2;
    T2[4351] = 2'h1;
    T2[4352] = 2'h2;
    T2[4353] = 2'h1;
    T2[4354] = 2'h3;
    T2[4355] = 2'h3;
    T2[4356] = 2'h1;
    T2[4357] = 2'h2;
    T2[4358] = 2'h1;
    T2[4359] = 2'h3;
    T2[4360] = 2'h0;
    T2[4361] = 2'h2;
    T2[4362] = 2'h2;
    T2[4363] = 2'h1;
    T2[4364] = 2'h3;
    T2[4365] = 2'h1;
    T2[4366] = 2'h2;
    T2[4367] = 2'h2;
    T2[4368] = 2'h1;
    T2[4369] = 2'h3;
    T2[4370] = 2'h2;
    T2[4371] = 2'h2;
    T2[4372] = 2'h2;
    T2[4373] = 2'h1;
    T2[4374] = 2'h3;
    T2[4375] = 2'h3;
    T2[4376] = 2'h2;
    T2[4377] = 2'h2;
    T2[4378] = 2'h1;
    T2[4379] = 2'h3;
    T2[4380] = 2'h0;
    T2[4381] = 2'h3;
    T2[4382] = 2'h2;
    T2[4383] = 2'h1;
    T2[4384] = 2'h3;
    T2[4385] = 2'h1;
    T2[4386] = 2'h3;
    T2[4387] = 2'h2;
    T2[4388] = 2'h1;
    T2[4389] = 2'h3;
    T2[4390] = 2'h2;
    T2[4391] = 2'h3;
    T2[4392] = 2'h2;
    T2[4393] = 2'h1;
    T2[4394] = 2'h3;
    T2[4395] = 2'h3;
    T2[4396] = 2'h3;
    T2[4397] = 2'h2;
    T2[4398] = 2'h1;
    T2[4399] = 2'h3;
    T2[4400] = 2'h0;
    T2[4401] = 2'h0;
    T2[4402] = 2'h3;
    T2[4403] = 2'h1;
    T2[4404] = 2'h3;
    T2[4405] = 2'h1;
    T2[4406] = 2'h0;
    T2[4407] = 2'h3;
    T2[4408] = 2'h1;
    T2[4409] = 2'h3;
    T2[4410] = 2'h2;
    T2[4411] = 2'h0;
    T2[4412] = 2'h3;
    T2[4413] = 2'h1;
    T2[4414] = 2'h3;
    T2[4415] = 2'h3;
    T2[4416] = 2'h0;
    T2[4417] = 2'h3;
    T2[4418] = 2'h1;
    T2[4419] = 2'h3;
    T2[4420] = 2'h0;
    T2[4421] = 2'h1;
    T2[4422] = 2'h3;
    T2[4423] = 2'h1;
    T2[4424] = 2'h3;
    T2[4425] = 2'h1;
    T2[4426] = 2'h1;
    T2[4427] = 2'h3;
    T2[4428] = 2'h1;
    T2[4429] = 2'h3;
    T2[4430] = 2'h2;
    T2[4431] = 2'h1;
    T2[4432] = 2'h3;
    T2[4433] = 2'h1;
    T2[4434] = 2'h3;
    T2[4435] = 2'h3;
    T2[4436] = 2'h1;
    T2[4437] = 2'h3;
    T2[4438] = 2'h1;
    T2[4439] = 2'h3;
    T2[4440] = 2'h0;
    T2[4441] = 2'h2;
    T2[4442] = 2'h3;
    T2[4443] = 2'h1;
    T2[4444] = 2'h3;
    T2[4445] = 2'h1;
    T2[4446] = 2'h2;
    T2[4447] = 2'h3;
    T2[4448] = 2'h1;
    T2[4449] = 2'h3;
    T2[4450] = 2'h2;
    T2[4451] = 2'h2;
    T2[4452] = 2'h3;
    T2[4453] = 2'h1;
    T2[4454] = 2'h3;
    T2[4455] = 2'h3;
    T2[4456] = 2'h2;
    T2[4457] = 2'h3;
    T2[4458] = 2'h1;
    T2[4459] = 2'h3;
    T2[4460] = 2'h0;
    T2[4461] = 2'h3;
    T2[4462] = 2'h3;
    T2[4463] = 2'h1;
    T2[4464] = 2'h3;
    T2[4465] = 2'h1;
    T2[4466] = 2'h3;
    T2[4467] = 2'h3;
    T2[4468] = 2'h1;
    T2[4469] = 2'h3;
    T2[4470] = 2'h2;
    T2[4471] = 2'h3;
    T2[4472] = 2'h3;
    T2[4473] = 2'h1;
    T2[4474] = 2'h3;
    T2[4475] = 2'h3;
    T2[4476] = 2'h3;
    T2[4477] = 2'h3;
    T2[4478] = 2'h1;
    T2[4479] = 2'h3;
    T2[4480] = 2'h0;
    T2[4481] = 2'h0;
    T2[4482] = 2'h0;
    T2[4483] = 2'h2;
    T2[4484] = 2'h3;
    T2[4485] = 2'h1;
    T2[4486] = 2'h0;
    T2[4487] = 2'h0;
    T2[4488] = 2'h2;
    T2[4489] = 2'h3;
    T2[4490] = 2'h2;
    T2[4491] = 2'h0;
    T2[4492] = 2'h0;
    T2[4493] = 2'h2;
    T2[4494] = 2'h3;
    T2[4495] = 2'h3;
    T2[4496] = 2'h0;
    T2[4497] = 2'h0;
    T2[4498] = 2'h2;
    T2[4499] = 2'h3;
    T2[4500] = 2'h0;
    T2[4501] = 2'h1;
    T2[4502] = 2'h0;
    T2[4503] = 2'h2;
    T2[4504] = 2'h3;
    T2[4505] = 2'h1;
    T2[4506] = 2'h1;
    T2[4507] = 2'h0;
    T2[4508] = 2'h2;
    T2[4509] = 2'h3;
    T2[4510] = 2'h2;
    T2[4511] = 2'h1;
    T2[4512] = 2'h0;
    T2[4513] = 2'h2;
    T2[4514] = 2'h3;
    T2[4515] = 2'h3;
    T2[4516] = 2'h1;
    T2[4517] = 2'h0;
    T2[4518] = 2'h2;
    T2[4519] = 2'h3;
    T2[4520] = 2'h0;
    T2[4521] = 2'h2;
    T2[4522] = 2'h0;
    T2[4523] = 2'h2;
    T2[4524] = 2'h3;
    T2[4525] = 2'h1;
    T2[4526] = 2'h2;
    T2[4527] = 2'h0;
    T2[4528] = 2'h2;
    T2[4529] = 2'h3;
    T2[4530] = 2'h2;
    T2[4531] = 2'h2;
    T2[4532] = 2'h0;
    T2[4533] = 2'h2;
    T2[4534] = 2'h3;
    T2[4535] = 2'h3;
    T2[4536] = 2'h2;
    T2[4537] = 2'h0;
    T2[4538] = 2'h2;
    T2[4539] = 2'h3;
    T2[4540] = 2'h0;
    T2[4541] = 2'h3;
    T2[4542] = 2'h0;
    T2[4543] = 2'h2;
    T2[4544] = 2'h3;
    T2[4545] = 2'h1;
    T2[4546] = 2'h3;
    T2[4547] = 2'h0;
    T2[4548] = 2'h2;
    T2[4549] = 2'h3;
    T2[4550] = 2'h2;
    T2[4551] = 2'h3;
    T2[4552] = 2'h0;
    T2[4553] = 2'h2;
    T2[4554] = 2'h3;
    T2[4555] = 2'h3;
    T2[4556] = 2'h3;
    T2[4557] = 2'h0;
    T2[4558] = 2'h2;
    T2[4559] = 2'h3;
    T2[4560] = 2'h0;
    T2[4561] = 2'h0;
    T2[4562] = 2'h1;
    T2[4563] = 2'h2;
    T2[4564] = 2'h3;
    T2[4565] = 2'h1;
    T2[4566] = 2'h0;
    T2[4567] = 2'h1;
    T2[4568] = 2'h2;
    T2[4569] = 2'h3;
    T2[4570] = 2'h2;
    T2[4571] = 2'h0;
    T2[4572] = 2'h1;
    T2[4573] = 2'h2;
    T2[4574] = 2'h3;
    T2[4575] = 2'h3;
    T2[4576] = 2'h0;
    T2[4577] = 2'h1;
    T2[4578] = 2'h2;
    T2[4579] = 2'h3;
    T2[4580] = 2'h0;
    T2[4581] = 2'h1;
    T2[4582] = 2'h1;
    T2[4583] = 2'h2;
    T2[4584] = 2'h3;
    T2[4585] = 2'h1;
    T2[4586] = 2'h1;
    T2[4587] = 2'h1;
    T2[4588] = 2'h2;
    T2[4589] = 2'h3;
    T2[4590] = 2'h2;
    T2[4591] = 2'h1;
    T2[4592] = 2'h1;
    T2[4593] = 2'h2;
    T2[4594] = 2'h3;
    T2[4595] = 2'h3;
    T2[4596] = 2'h1;
    T2[4597] = 2'h1;
    T2[4598] = 2'h2;
    T2[4599] = 2'h3;
    T2[4600] = 2'h0;
    T2[4601] = 2'h2;
    T2[4602] = 2'h1;
    T2[4603] = 2'h2;
    T2[4604] = 2'h3;
    T2[4605] = 2'h1;
    T2[4606] = 2'h2;
    T2[4607] = 2'h1;
    T2[4608] = 2'h2;
    T2[4609] = 2'h3;
    T2[4610] = 2'h2;
    T2[4611] = 2'h2;
    T2[4612] = 2'h1;
    T2[4613] = 2'h2;
    T2[4614] = 2'h3;
    T2[4615] = 2'h3;
    T2[4616] = 2'h2;
    T2[4617] = 2'h1;
    T2[4618] = 2'h2;
    T2[4619] = 2'h3;
    T2[4620] = 2'h0;
    T2[4621] = 2'h3;
    T2[4622] = 2'h1;
    T2[4623] = 2'h2;
    T2[4624] = 2'h3;
    T2[4625] = 2'h1;
    T2[4626] = 2'h3;
    T2[4627] = 2'h1;
    T2[4628] = 2'h2;
    T2[4629] = 2'h3;
    T2[4630] = 2'h2;
    T2[4631] = 2'h3;
    T2[4632] = 2'h1;
    T2[4633] = 2'h2;
    T2[4634] = 2'h3;
    T2[4635] = 2'h3;
    T2[4636] = 2'h3;
    T2[4637] = 2'h1;
    T2[4638] = 2'h2;
    T2[4639] = 2'h3;
    T2[4640] = 2'h0;
    T2[4641] = 2'h0;
    T2[4642] = 2'h2;
    T2[4643] = 2'h2;
    T2[4644] = 2'h3;
    T2[4645] = 2'h1;
    T2[4646] = 2'h0;
    T2[4647] = 2'h2;
    T2[4648] = 2'h2;
    T2[4649] = 2'h3;
    T2[4650] = 2'h2;
    T2[4651] = 2'h0;
    T2[4652] = 2'h2;
    T2[4653] = 2'h2;
    T2[4654] = 2'h3;
    T2[4655] = 2'h3;
    T2[4656] = 2'h0;
    T2[4657] = 2'h2;
    T2[4658] = 2'h2;
    T2[4659] = 2'h3;
    T2[4660] = 2'h0;
    T2[4661] = 2'h1;
    T2[4662] = 2'h2;
    T2[4663] = 2'h2;
    T2[4664] = 2'h3;
    T2[4665] = 2'h1;
    T2[4666] = 2'h1;
    T2[4667] = 2'h2;
    T2[4668] = 2'h2;
    T2[4669] = 2'h3;
    T2[4670] = 2'h2;
    T2[4671] = 2'h1;
    T2[4672] = 2'h2;
    T2[4673] = 2'h2;
    T2[4674] = 2'h3;
    T2[4675] = 2'h3;
    T2[4676] = 2'h1;
    T2[4677] = 2'h2;
    T2[4678] = 2'h2;
    T2[4679] = 2'h3;
    T2[4680] = 2'h0;
    T2[4681] = 2'h2;
    T2[4682] = 2'h2;
    T2[4683] = 2'h2;
    T2[4684] = 2'h3;
    T2[4685] = 2'h1;
    T2[4686] = 2'h2;
    T2[4687] = 2'h2;
    T2[4688] = 2'h2;
    T2[4689] = 2'h3;
    T2[4690] = 2'h2;
    T2[4691] = 2'h2;
    T2[4692] = 2'h2;
    T2[4693] = 2'h2;
    T2[4694] = 2'h3;
    T2[4695] = 2'h3;
    T2[4696] = 2'h2;
    T2[4697] = 2'h2;
    T2[4698] = 2'h2;
    T2[4699] = 2'h3;
    T2[4700] = 2'h0;
    T2[4701] = 2'h3;
    T2[4702] = 2'h2;
    T2[4703] = 2'h2;
    T2[4704] = 2'h3;
    T2[4705] = 2'h1;
    T2[4706] = 2'h3;
    T2[4707] = 2'h2;
    T2[4708] = 2'h2;
    T2[4709] = 2'h3;
    T2[4710] = 2'h2;
    T2[4711] = 2'h3;
    T2[4712] = 2'h2;
    T2[4713] = 2'h2;
    T2[4714] = 2'h3;
    T2[4715] = 2'h3;
    T2[4716] = 2'h3;
    T2[4717] = 2'h2;
    T2[4718] = 2'h2;
    T2[4719] = 2'h3;
    T2[4720] = 2'h0;
    T2[4721] = 2'h0;
    T2[4722] = 2'h3;
    T2[4723] = 2'h2;
    T2[4724] = 2'h3;
    T2[4725] = 2'h1;
    T2[4726] = 2'h0;
    T2[4727] = 2'h3;
    T2[4728] = 2'h2;
    T2[4729] = 2'h3;
    T2[4730] = 2'h2;
    T2[4731] = 2'h0;
    T2[4732] = 2'h3;
    T2[4733] = 2'h2;
    T2[4734] = 2'h3;
    T2[4735] = 2'h3;
    T2[4736] = 2'h0;
    T2[4737] = 2'h3;
    T2[4738] = 2'h2;
    T2[4739] = 2'h3;
    T2[4740] = 2'h0;
    T2[4741] = 2'h1;
    T2[4742] = 2'h3;
    T2[4743] = 2'h2;
    T2[4744] = 2'h3;
    T2[4745] = 2'h1;
    T2[4746] = 2'h1;
    T2[4747] = 2'h3;
    T2[4748] = 2'h2;
    T2[4749] = 2'h3;
    T2[4750] = 2'h2;
    T2[4751] = 2'h1;
    T2[4752] = 2'h3;
    T2[4753] = 2'h2;
    T2[4754] = 2'h3;
    T2[4755] = 2'h3;
    T2[4756] = 2'h1;
    T2[4757] = 2'h3;
    T2[4758] = 2'h2;
    T2[4759] = 2'h3;
    T2[4760] = 2'h0;
    T2[4761] = 2'h2;
    T2[4762] = 2'h3;
    T2[4763] = 2'h2;
    T2[4764] = 2'h3;
    T2[4765] = 2'h1;
    T2[4766] = 2'h2;
    T2[4767] = 2'h3;
    T2[4768] = 2'h2;
    T2[4769] = 2'h3;
    T2[4770] = 2'h2;
    T2[4771] = 2'h2;
    T2[4772] = 2'h3;
    T2[4773] = 2'h2;
    T2[4774] = 2'h3;
    T2[4775] = 2'h3;
    T2[4776] = 2'h2;
    T2[4777] = 2'h3;
    T2[4778] = 2'h2;
    T2[4779] = 2'h3;
    T2[4780] = 2'h0;
    T2[4781] = 2'h3;
    T2[4782] = 2'h3;
    T2[4783] = 2'h2;
    T2[4784] = 2'h3;
    T2[4785] = 2'h1;
    T2[4786] = 2'h3;
    T2[4787] = 2'h3;
    T2[4788] = 2'h2;
    T2[4789] = 2'h3;
    T2[4790] = 2'h2;
    T2[4791] = 2'h3;
    T2[4792] = 2'h3;
    T2[4793] = 2'h2;
    T2[4794] = 2'h3;
    T2[4795] = 2'h3;
    T2[4796] = 2'h3;
    T2[4797] = 2'h3;
    T2[4798] = 2'h2;
    T2[4799] = 2'h3;
    T2[4800] = 2'h0;
    T2[4801] = 2'h0;
    T2[4802] = 2'h0;
    T2[4803] = 2'h3;
    T2[4804] = 2'h3;
    T2[4805] = 2'h1;
    T2[4806] = 2'h0;
    T2[4807] = 2'h0;
    T2[4808] = 2'h3;
    T2[4809] = 2'h3;
    T2[4810] = 2'h2;
    T2[4811] = 2'h0;
    T2[4812] = 2'h0;
    T2[4813] = 2'h3;
    T2[4814] = 2'h3;
    T2[4815] = 2'h3;
    T2[4816] = 2'h0;
    T2[4817] = 2'h0;
    T2[4818] = 2'h3;
    T2[4819] = 2'h3;
    T2[4820] = 2'h0;
    T2[4821] = 2'h1;
    T2[4822] = 2'h0;
    T2[4823] = 2'h3;
    T2[4824] = 2'h3;
    T2[4825] = 2'h1;
    T2[4826] = 2'h1;
    T2[4827] = 2'h0;
    T2[4828] = 2'h3;
    T2[4829] = 2'h3;
    T2[4830] = 2'h2;
    T2[4831] = 2'h1;
    T2[4832] = 2'h0;
    T2[4833] = 2'h3;
    T2[4834] = 2'h3;
    T2[4835] = 2'h3;
    T2[4836] = 2'h1;
    T2[4837] = 2'h0;
    T2[4838] = 2'h3;
    T2[4839] = 2'h3;
    T2[4840] = 2'h0;
    T2[4841] = 2'h2;
    T2[4842] = 2'h0;
    T2[4843] = 2'h3;
    T2[4844] = 2'h3;
    T2[4845] = 2'h1;
    T2[4846] = 2'h2;
    T2[4847] = 2'h0;
    T2[4848] = 2'h3;
    T2[4849] = 2'h3;
    T2[4850] = 2'h2;
    T2[4851] = 2'h2;
    T2[4852] = 2'h0;
    T2[4853] = 2'h3;
    T2[4854] = 2'h3;
    T2[4855] = 2'h3;
    T2[4856] = 2'h2;
    T2[4857] = 2'h0;
    T2[4858] = 2'h3;
    T2[4859] = 2'h3;
    T2[4860] = 2'h0;
    T2[4861] = 2'h3;
    T2[4862] = 2'h0;
    T2[4863] = 2'h3;
    T2[4864] = 2'h3;
    T2[4865] = 2'h1;
    T2[4866] = 2'h3;
    T2[4867] = 2'h0;
    T2[4868] = 2'h3;
    T2[4869] = 2'h3;
    T2[4870] = 2'h2;
    T2[4871] = 2'h3;
    T2[4872] = 2'h0;
    T2[4873] = 2'h3;
    T2[4874] = 2'h3;
    T2[4875] = 2'h3;
    T2[4876] = 2'h3;
    T2[4877] = 2'h0;
    T2[4878] = 2'h3;
    T2[4879] = 2'h3;
    T2[4880] = 2'h0;
    T2[4881] = 2'h0;
    T2[4882] = 2'h1;
    T2[4883] = 2'h3;
    T2[4884] = 2'h3;
    T2[4885] = 2'h1;
    T2[4886] = 2'h0;
    T2[4887] = 2'h1;
    T2[4888] = 2'h3;
    T2[4889] = 2'h3;
    T2[4890] = 2'h2;
    T2[4891] = 2'h0;
    T2[4892] = 2'h1;
    T2[4893] = 2'h3;
    T2[4894] = 2'h3;
    T2[4895] = 2'h3;
    T2[4896] = 2'h0;
    T2[4897] = 2'h1;
    T2[4898] = 2'h3;
    T2[4899] = 2'h3;
    T2[4900] = 2'h0;
    T2[4901] = 2'h1;
    T2[4902] = 2'h1;
    T2[4903] = 2'h3;
    T2[4904] = 2'h3;
    T2[4905] = 2'h1;
    T2[4906] = 2'h1;
    T2[4907] = 2'h1;
    T2[4908] = 2'h3;
    T2[4909] = 2'h3;
    T2[4910] = 2'h2;
    T2[4911] = 2'h1;
    T2[4912] = 2'h1;
    T2[4913] = 2'h3;
    T2[4914] = 2'h3;
    T2[4915] = 2'h3;
    T2[4916] = 2'h1;
    T2[4917] = 2'h1;
    T2[4918] = 2'h3;
    T2[4919] = 2'h3;
    T2[4920] = 2'h0;
    T2[4921] = 2'h2;
    T2[4922] = 2'h1;
    T2[4923] = 2'h3;
    T2[4924] = 2'h3;
    T2[4925] = 2'h1;
    T2[4926] = 2'h2;
    T2[4927] = 2'h1;
    T2[4928] = 2'h3;
    T2[4929] = 2'h3;
    T2[4930] = 2'h2;
    T2[4931] = 2'h2;
    T2[4932] = 2'h1;
    T2[4933] = 2'h3;
    T2[4934] = 2'h3;
    T2[4935] = 2'h3;
    T2[4936] = 2'h2;
    T2[4937] = 2'h1;
    T2[4938] = 2'h3;
    T2[4939] = 2'h3;
    T2[4940] = 2'h0;
    T2[4941] = 2'h3;
    T2[4942] = 2'h1;
    T2[4943] = 2'h3;
    T2[4944] = 2'h3;
    T2[4945] = 2'h1;
    T2[4946] = 2'h3;
    T2[4947] = 2'h1;
    T2[4948] = 2'h3;
    T2[4949] = 2'h3;
    T2[4950] = 2'h2;
    T2[4951] = 2'h3;
    T2[4952] = 2'h1;
    T2[4953] = 2'h3;
    T2[4954] = 2'h3;
    T2[4955] = 2'h3;
    T2[4956] = 2'h3;
    T2[4957] = 2'h1;
    T2[4958] = 2'h3;
    T2[4959] = 2'h3;
    T2[4960] = 2'h0;
    T2[4961] = 2'h0;
    T2[4962] = 2'h2;
    T2[4963] = 2'h3;
    T2[4964] = 2'h3;
    T2[4965] = 2'h1;
    T2[4966] = 2'h0;
    T2[4967] = 2'h2;
    T2[4968] = 2'h3;
    T2[4969] = 2'h3;
    T2[4970] = 2'h2;
    T2[4971] = 2'h0;
    T2[4972] = 2'h2;
    T2[4973] = 2'h3;
    T2[4974] = 2'h3;
    T2[4975] = 2'h3;
    T2[4976] = 2'h0;
    T2[4977] = 2'h2;
    T2[4978] = 2'h3;
    T2[4979] = 2'h3;
    T2[4980] = 2'h0;
    T2[4981] = 2'h1;
    T2[4982] = 2'h2;
    T2[4983] = 2'h3;
    T2[4984] = 2'h3;
    T2[4985] = 2'h1;
    T2[4986] = 2'h1;
    T2[4987] = 2'h2;
    T2[4988] = 2'h3;
    T2[4989] = 2'h3;
    T2[4990] = 2'h2;
    T2[4991] = 2'h1;
    T2[4992] = 2'h2;
    T2[4993] = 2'h3;
    T2[4994] = 2'h3;
    T2[4995] = 2'h3;
    T2[4996] = 2'h1;
    T2[4997] = 2'h2;
    T2[4998] = 2'h3;
    T2[4999] = 2'h3;
    T2[5000] = 2'h0;
    T2[5001] = 2'h2;
    T2[5002] = 2'h2;
    T2[5003] = 2'h3;
    T2[5004] = 2'h3;
    T2[5005] = 2'h1;
    T2[5006] = 2'h2;
    T2[5007] = 2'h2;
    T2[5008] = 2'h3;
    T2[5009] = 2'h3;
    T2[5010] = 2'h2;
    T2[5011] = 2'h2;
    T2[5012] = 2'h2;
    T2[5013] = 2'h3;
    T2[5014] = 2'h3;
    T2[5015] = 2'h3;
    T2[5016] = 2'h2;
    T2[5017] = 2'h2;
    T2[5018] = 2'h3;
    T2[5019] = 2'h3;
    T2[5020] = 2'h0;
    T2[5021] = 2'h3;
    T2[5022] = 2'h2;
    T2[5023] = 2'h3;
    T2[5024] = 2'h3;
    T2[5025] = 2'h1;
    T2[5026] = 2'h3;
    T2[5027] = 2'h2;
    T2[5028] = 2'h3;
    T2[5029] = 2'h3;
    T2[5030] = 2'h2;
    T2[5031] = 2'h3;
    T2[5032] = 2'h2;
    T2[5033] = 2'h3;
    T2[5034] = 2'h3;
    T2[5035] = 2'h3;
    T2[5036] = 2'h3;
    T2[5037] = 2'h2;
    T2[5038] = 2'h3;
    T2[5039] = 2'h3;
    T2[5040] = 2'h0;
    T2[5041] = 2'h0;
    T2[5042] = 2'h3;
    T2[5043] = 2'h3;
    T2[5044] = 2'h3;
    T2[5045] = 2'h1;
    T2[5046] = 2'h0;
    T2[5047] = 2'h3;
    T2[5048] = 2'h3;
    T2[5049] = 2'h3;
    T2[5050] = 2'h2;
    T2[5051] = 2'h0;
    T2[5052] = 2'h3;
    T2[5053] = 2'h3;
    T2[5054] = 2'h3;
    T2[5055] = 2'h3;
    T2[5056] = 2'h0;
    T2[5057] = 2'h3;
    T2[5058] = 2'h3;
    T2[5059] = 2'h3;
    T2[5060] = 2'h0;
    T2[5061] = 2'h1;
    T2[5062] = 2'h3;
    T2[5063] = 2'h3;
    T2[5064] = 2'h3;
    T2[5065] = 2'h1;
    T2[5066] = 2'h1;
    T2[5067] = 2'h3;
    T2[5068] = 2'h3;
    T2[5069] = 2'h3;
    T2[5070] = 2'h2;
    T2[5071] = 2'h1;
    T2[5072] = 2'h3;
    T2[5073] = 2'h3;
    T2[5074] = 2'h3;
    T2[5075] = 2'h3;
    T2[5076] = 2'h1;
    T2[5077] = 2'h3;
    T2[5078] = 2'h3;
    T2[5079] = 2'h3;
    T2[5080] = 2'h0;
    T2[5081] = 2'h2;
    T2[5082] = 2'h3;
    T2[5083] = 2'h3;
    T2[5084] = 2'h3;
    T2[5085] = 2'h1;
    T2[5086] = 2'h2;
    T2[5087] = 2'h3;
    T2[5088] = 2'h3;
    T2[5089] = 2'h3;
    T2[5090] = 2'h2;
    T2[5091] = 2'h2;
    T2[5092] = 2'h3;
    T2[5093] = 2'h3;
    T2[5094] = 2'h3;
    T2[5095] = 2'h3;
    T2[5096] = 2'h2;
    T2[5097] = 2'h3;
    T2[5098] = 2'h3;
    T2[5099] = 2'h3;
    T2[5100] = 2'h0;
    T2[5101] = 2'h3;
    T2[5102] = 2'h3;
    T2[5103] = 2'h3;
    T2[5104] = 2'h3;
    T2[5105] = 2'h1;
    T2[5106] = 2'h3;
    T2[5107] = 2'h3;
    T2[5108] = 2'h3;
    T2[5109] = 2'h3;
    T2[5110] = 2'h2;
    T2[5111] = 2'h3;
    T2[5112] = 2'h3;
    T2[5113] = 2'h3;
    T2[5114] = 2'h3;
    T2[5115] = 2'h3;
    T2[5116] = 2'h3;
    T2[5117] = 2'h3;
    T2[5118] = 2'h3;
    T2[5119] = 2'h3;
  end
  assign T3 = T4[4'hc:1'h0];
  assign T4 = index + T5;
  assign T5 = {11'h0, io_inb};
  assign index = io_ina * 3'h5;
endmodule

