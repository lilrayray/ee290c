module powerLUT(
    input [5:0] io_fftsize,
    input [2:0] io_power,
    output[2:0] io_power4235
);

  wire[2:0] T0;
  reg [2:0] T1 [167:0];
  wire[7:0] T2;


  assign io_power4235 = T0;
`ifndef SYNTHESIS
  assign T0 = T2 >= 8'ha8 ? {1{$random}} : T1[T2];
`else
  assign T0 = T1[T2];
`endif
  always @(*) begin
    T1[0] = 3'h1;
    T1[1] = 3'h0;
    T1[2] = 3'h1;
    T1[3] = 3'h0;
    T1[4] = 3'h1;
    T1[5] = 3'h1;
    T1[6] = 3'h1;
    T1[7] = 3'h0;
    T1[8] = 3'h1;
    T1[9] = 3'h0;
    T1[10] = 3'h2;
    T1[11] = 3'h0;
    T1[12] = 3'h2;
    T1[13] = 3'h0;
    T1[14] = 3'h1;
    T1[15] = 3'h0;
    T1[16] = 3'h1;
    T1[17] = 3'h0;
    T1[18] = 3'h1;
    T1[19] = 3'h1;
    T1[20] = 3'h1;
    T1[21] = 3'h1;
    T1[22] = 3'h2;
    T1[23] = 3'h0;
    T1[24] = 3'h2;
    T1[25] = 3'h1;
    T1[26] = 3'h1;
    T1[27] = 3'h0;
    T1[28] = 3'h1;
    T1[29] = 3'h0;
    T1[30] = 3'h3;
    T1[31] = 3'h0;
    T1[32] = 3'h1;
    T1[33] = 3'h1;
    T1[34] = 3'h1;
    T1[35] = 3'h1;
    T1[36] = 3'h2;
    T1[37] = 3'h0;
    T1[38] = 3'h2;
    T1[39] = 3'h0;
    T1[40] = 3'h1;
    T1[41] = 3'h0;
    T1[42] = 3'h2;
    T1[43] = 3'h1;
    T1[44] = 3'h3;
    T1[45] = 3'h0;
    T1[46] = 3'h1;
    T1[47] = 3'h0;
    T1[48] = 3'h1;
    T1[49] = 3'h1;
    T1[50] = 3'h3;
    T1[51] = 3'h0;
    T1[52] = 3'h2;
    T1[53] = 3'h0;
    T1[54] = 3'h1;
    T1[55] = 3'h1;
    T1[56] = 3'h2;
    T1[57] = 3'h1;
    T1[58] = 3'h2;
    T1[59] = 3'h0;
    T1[60] = 3'h1;
    T1[61] = 3'h0;
    T1[62] = 3'h1;
    T1[63] = 3'h2;
    T1[64] = 3'h1;
    T1[65] = 3'h0;
    T1[66] = 3'h4;
    T1[67] = 3'h0;
    T1[68] = 3'h1;
    T1[69] = 3'h1;
    T1[70] = 3'h2;
    T1[71] = 3'h1;
    T1[72] = 3'h3;
    T1[73] = 3'h1;
    T1[74] = 3'h1;
    T1[75] = 3'h0;
    T1[76] = 3'h2;
    T1[77] = 3'h0;
    T1[78] = 3'h3;
    T1[79] = 3'h0;
    T1[80] = 3'h2;
    T1[81] = 3'h1;
    T1[82] = 3'h1;
    T1[83] = 3'h1;
    T1[84] = 3'h1;
    T1[85] = 3'h0;
    T1[86] = 3'h3;
    T1[87] = 3'h1;
    T1[88] = 3'h3;
    T1[89] = 3'h0;
    T1[90] = 3'h2;
    T1[91] = 3'h0;
    T1[92] = 3'h1;
    T1[93] = 3'h1;
    T1[94] = 3'h1;
    T1[95] = 3'h2;
    T1[96] = 3'h1;
    T1[97] = 3'h1;
    T1[98] = 3'h4;
    T1[99] = 3'h0;
    T1[100] = 3'h2;
    T1[101] = 3'h0;
    T1[102] = 3'h2;
    T1[103] = 3'h1;
    T1[104] = 3'h4;
    T1[105] = 3'h0;
    T1[106] = 3'h1;
    T1[107] = 3'h0;
    T1[108] = 3'h2;
    T1[109] = 3'h1;
    T1[110] = 3'h3;
    T1[111] = 3'h0;
    T1[112] = 3'h1;
    T1[113] = 3'h0;
    T1[114] = 3'h2;
    T1[115] = 3'h2;
    T1[116] = 3'h3;
    T1[117] = 3'h0;
    T1[118] = 3'h1;
    T1[119] = 3'h1;
    T1[120] = 3'h1;
    T1[121] = 3'h0;
    T1[122] = 3'h5;
    T1[123] = 3'h0;
    T1[124] = 3'h1;
    T1[125] = 3'h1;
    T1[126] = 3'h3;
    T1[127] = 3'h1;
    T1[128] = 3'h3;
    T1[129] = 3'h1;
    T1[130] = 3'h2;
    T1[131] = 3'h0;
    T1[132] = 3'h2;
    T1[133] = 3'h0;
    T1[134] = 3'h1;
    T1[135] = 3'h2;
    T1[136] = 3'h2;
    T1[137] = 3'h0;
    T1[138] = 3'h4;
    T1[139] = 3'h0;
    T1[140] = 3'h4;
    T1[141] = 3'h1;
    T1[142] = 3'h1;
    T1[143] = 3'h0;
    T1[144] = 3'h3;
    T1[145] = 3'h0;
    T1[146] = 3'h0;
    T1[147] = 3'h0;
    T1[148] = 3'h3;
    T1[149] = 3'h1;
    T1[150] = 3'h0;
    T1[151] = 3'h0;
    T1[152] = 3'h4;
    T1[153] = 3'h0;
    T1[154] = 3'h0;
    T1[155] = 3'h0;
    T1[156] = 3'h4;
    T1[157] = 3'h1;
    T1[158] = 3'h0;
    T1[159] = 3'h0;
    T1[160] = 3'h5;
    T1[161] = 3'h0;
    T1[162] = 3'h0;
    T1[163] = 3'h0;
    T1[164] = 3'h5;
    T1[165] = 3'h1;
    T1[166] = 3'h0;
    T1[167] = 3'h0;
  end
  assign T2 = {2'h0, io_fftsize};
endmodule

