module twiddleLUT(
    input [9:0] io_in4,
    input [9:0] io_in5,
    input [9:0] io_in3,
    output[15:0] io_t4_1out_real,
    output[15:0] io_t4_1out_imag,
    output[15:0] io_t4_2out_real,
    output[15:0] io_t4_2out_imag,
    output[15:0] io_t4_3out_real,
    output[15:0] io_t4_3out_imag,
    output[15:0] io_t3_1out_real,
    output[15:0] io_t3_1out_imag,
    output[15:0] io_t3_2out_real,
    output[15:0] io_t3_2out_imag,
    output[15:0] io_t5_1out_real,
    output[15:0] io_t5_1out_imag,
    output[15:0] io_t5_2out_real,
    output[15:0] io_t5_2out_imag,
    output[15:0] io_t5_3out_real,
    output[15:0] io_t5_3out_imag,
    output[15:0] io_t5_4out_real,
    output[15:0] io_t5_4out_imag
);

  wire[15:0] T0;
  wire[47:0] T1;
  wire[47:0] T2;
  wire[47:0] T3;
  wire[47:0] twiddle5_4_0_imag;
  wire[47:0] T4;
  wire[16:0] T5;
  wire[16:0] T6;
  wire[30:0] T7;
  wire T8;
  wire[47:0] T9;
  wire[47:0] T10;
  wire[47:0] T11;
  wire[46:0] twiddle5_4_1_imag;
  wire[46:0] T12;
  wire[46:0] T13;
  wire[46:0] T14;
  wire[46:0] T15;
  wire T16;
  wire T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[47:0] T20;
  wire[46:0] T21;
  wire[46:0] twiddle5_4_2_imag;
  wire[46:0] T22;
  wire[46:0] T23;
  wire[46:0] T24;
  wire[45:0] T25;
  wire[45:0] T26;
  wire T27;
  wire[46:0] twiddle5_4_3_imag;
  wire[46:0] T28;
  wire[44:0] T29;
  wire[44:0] T30;
  wire[1:0] T31;
  wire T32;
  wire[46:0] T33;
  wire[46:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire[47:0] T38;
  wire[46:0] twiddle5_4_4_imag;
  wire[46:0] T39;
  wire[46:0] T40;
  wire[46:0] T41;
  wire[46:0] T42;
  wire T43;
  wire T44;
  wire[15:0] T45;
  wire[47:0] T46;
  wire[47:0] T47;
  wire[47:0] T48;
  wire[47:0] twiddle5_4_0_real;
  wire[47:0] T49;
  wire[16:0] T50;
  wire[16:0] T51;
  wire[30:0] T52;
  wire T53;
  wire[47:0] T54;
  wire[47:0] T55;
  wire[47:0] T56;
  wire[46:0] twiddle5_4_1_real;
  wire[46:0] T57;
  wire[46:0] T58;
  wire[46:0] T59;
  wire[46:0] T60;
  wire T61;
  wire T62;
  wire[47:0] T63;
  wire[46:0] T64;
  wire[46:0] twiddle5_4_2_real;
  wire[46:0] T65;
  wire[46:0] T66;
  wire[46:0] T67;
  wire[45:0] T68;
  wire[45:0] T69;
  wire T70;
  wire[46:0] twiddle5_4_3_real;
  wire[46:0] T71;
  wire[44:0] T72;
  wire[44:0] T73;
  wire[1:0] T74;
  wire T75;
  wire[46:0] T76;
  wire[46:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[47:0] T81;
  wire[46:0] twiddle5_4_4_real;
  wire[46:0] T82;
  wire[46:0] T83;
  wire[46:0] T84;
  wire[46:0] T85;
  wire T86;
  wire T87;
  wire[15:0] T88;
  wire[47:0] T89;
  wire[47:0] T90;
  wire[47:0] T91;
  wire[47:0] twiddle5_3_0_imag;
  wire[47:0] T92;
  wire[16:0] T93;
  wire[16:0] T94;
  wire[30:0] T95;
  wire T96;
  wire[47:0] T97;
  wire[47:0] T98;
  wire[47:0] T99;
  wire[46:0] twiddle5_3_1_imag;
  wire[46:0] T100;
  wire[46:0] T101;
  wire[46:0] T102;
  wire[46:0] T103;
  wire T104;
  wire T105;
  wire[2:0] T106;
  wire[2:0] T107;
  wire[47:0] T108;
  wire[46:0] T109;
  wire[46:0] twiddle5_3_2_imag;
  wire[46:0] T110;
  wire[46:0] T111;
  wire[46:0] T112;
  wire[43:0] T113;
  wire[43:0] T114;
  wire[2:0] T115;
  wire T116;
  wire[46:0] twiddle5_3_3_imag;
  wire[46:0] T117;
  wire[46:0] T118;
  wire[46:0] T119;
  wire[46:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire[47:0] T124;
  wire[46:0] twiddle5_3_4_imag;
  wire[46:0] T125;
  wire[44:0] T126;
  wire[44:0] T127;
  wire[1:0] T128;
  wire T129;
  wire[46:0] T130;
  wire[46:0] T131;
  wire T132;
  wire T133;
  wire[15:0] T134;
  wire[47:0] T135;
  wire[47:0] T136;
  wire[47:0] T137;
  wire[47:0] twiddle5_3_0_real;
  wire[47:0] T138;
  wire[16:0] T139;
  wire[16:0] T140;
  wire[30:0] T141;
  wire T142;
  wire[47:0] T143;
  wire[47:0] T144;
  wire[47:0] T145;
  wire[46:0] twiddle5_3_1_real;
  wire[46:0] T146;
  wire[46:0] T147;
  wire[46:0] T148;
  wire[46:0] T149;
  wire T150;
  wire T151;
  wire[47:0] T152;
  wire[46:0] T153;
  wire[46:0] twiddle5_3_2_real;
  wire[46:0] T154;
  wire[46:0] T155;
  wire[46:0] T156;
  wire[43:0] T157;
  wire[43:0] T158;
  wire[2:0] T159;
  wire T160;
  wire[46:0] twiddle5_3_3_real;
  wire[46:0] T161;
  wire[46:0] T162;
  wire[46:0] T163;
  wire[46:0] T164;
  wire T165;
  wire T166;
  wire T167;
  wire[47:0] T168;
  wire[46:0] twiddle5_3_4_real;
  wire[46:0] T169;
  wire[44:0] T170;
  wire[44:0] T171;
  wire[1:0] T172;
  wire T173;
  wire[46:0] T174;
  wire[46:0] T175;
  wire T176;
  wire T177;
  wire[15:0] T178;
  wire[47:0] T179;
  wire[47:0] T180;
  wire[47:0] T181;
  wire[47:0] twiddle5_2_0_imag;
  wire[47:0] T182;
  wire[16:0] T183;
  wire[16:0] T184;
  wire[30:0] T185;
  wire T186;
  wire[47:0] T187;
  wire[47:0] T188;
  wire[47:0] T189;
  wire[46:0] twiddle5_2_1_imag;
  wire[46:0] T190;
  wire[45:0] T191;
  wire[45:0] T192;
  wire T193;
  wire[46:0] T194;
  wire[46:0] T195;
  wire T196;
  wire T197;
  wire[2:0] T198;
  wire[2:0] T199;
  wire[47:0] T200;
  wire[46:0] T201;
  wire[46:0] twiddle5_2_2_imag;
  wire[46:0] T202;
  wire[46:0] T203;
  wire[46:0] T204;
  wire[46:0] T205;
  wire[46:0] twiddle5_2_3_imag;
  wire[46:0] T206;
  wire[46:0] T207;
  wire[46:0] T208;
  wire[43:0] T209;
  wire[43:0] T210;
  wire[2:0] T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire[47:0] T216;
  wire[46:0] twiddle5_2_4_imag;
  wire[46:0] T217;
  wire[46:0] T218;
  wire[46:0] T219;
  wire[45:0] T220;
  wire[45:0] T221;
  wire T222;
  wire T223;
  wire T224;
  wire[15:0] T225;
  wire[47:0] T226;
  wire[47:0] T227;
  wire[47:0] T228;
  wire[47:0] twiddle5_2_0_real;
  wire[47:0] T229;
  wire[16:0] T230;
  wire[16:0] T231;
  wire[30:0] T232;
  wire T233;
  wire[47:0] T234;
  wire[47:0] T235;
  wire[47:0] T236;
  wire[46:0] twiddle5_2_1_real;
  wire[46:0] T237;
  wire[45:0] T238;
  wire[45:0] T239;
  wire T240;
  wire[46:0] T241;
  wire[46:0] T242;
  wire T243;
  wire T244;
  wire[47:0] T245;
  wire[46:0] T246;
  wire[46:0] twiddle5_2_2_real;
  wire[46:0] T247;
  wire[46:0] T248;
  wire[46:0] T249;
  wire[46:0] T250;
  wire[46:0] twiddle5_2_3_real;
  wire[46:0] T251;
  wire[46:0] T252;
  wire[46:0] T253;
  wire[43:0] T254;
  wire[43:0] T255;
  wire[2:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire[47:0] T261;
  wire[46:0] twiddle5_2_4_real;
  wire[46:0] T262;
  wire[46:0] T263;
  wire[46:0] T264;
  wire[45:0] T265;
  wire[45:0] T266;
  wire T267;
  wire T268;
  wire T269;
  wire[15:0] T270;
  wire[47:0] T271;
  wire[47:0] T272;
  wire[47:0] T273;
  wire[47:0] twiddle5_1_0_imag;
  wire[47:0] T274;
  wire[16:0] T275;
  wire[16:0] T276;
  wire[30:0] T277;
  wire T278;
  wire[47:0] T279;
  wire[47:0] T280;
  wire[47:0] T281;
  wire[46:0] twiddle5_1_1_imag;
  wire[46:0] T282;
  wire[44:0] T283;
  wire[44:0] T284;
  wire[1:0] T285;
  wire T286;
  wire[46:0] T287;
  wire[46:0] T288;
  wire T289;
  wire T290;
  wire[2:0] T291;
  wire[2:0] T292;
  wire[47:0] T293;
  wire[46:0] T294;
  wire[46:0] twiddle5_1_2_imag;
  wire[46:0] T295;
  wire[45:0] T296;
  wire[45:0] T297;
  wire T298;
  wire[46:0] T299;
  wire[46:0] T300;
  wire[46:0] twiddle5_1_3_imag;
  wire[46:0] T301;
  wire[46:0] T302;
  wire[46:0] T303;
  wire[46:0] T304;
  wire T305;
  wire T306;
  wire T307;
  wire[47:0] T308;
  wire[46:0] twiddle5_1_4_imag;
  wire[46:0] T309;
  wire[46:0] T310;
  wire[46:0] T311;
  wire[46:0] T312;
  wire T313;
  wire T314;
  wire[15:0] T315;
  wire[47:0] T316;
  wire[47:0] T317;
  wire[47:0] T318;
  wire[47:0] twiddle5_1_0_real;
  wire[47:0] T319;
  wire[16:0] T320;
  wire[16:0] T321;
  wire[30:0] T322;
  wire T323;
  wire[47:0] T324;
  wire[47:0] T325;
  wire[47:0] T326;
  wire[46:0] twiddle5_1_1_real;
  wire[46:0] T327;
  wire[44:0] T328;
  wire[44:0] T329;
  wire[1:0] T330;
  wire T331;
  wire[46:0] T332;
  wire[46:0] T333;
  wire T334;
  wire T335;
  wire[47:0] T336;
  wire[46:0] T337;
  wire[46:0] twiddle5_1_2_real;
  wire[46:0] T338;
  wire[45:0] T339;
  wire[45:0] T340;
  wire T341;
  wire[46:0] T342;
  wire[46:0] T343;
  wire[46:0] twiddle5_1_3_real;
  wire[46:0] T344;
  wire[46:0] T345;
  wire[46:0] T346;
  wire[46:0] T347;
  wire T348;
  wire T349;
  wire T350;
  wire[47:0] T351;
  wire[46:0] twiddle5_1_4_real;
  wire[46:0] T352;
  wire[46:0] T353;
  wire[46:0] T354;
  wire[46:0] T355;
  wire T356;
  wire T357;
  wire[15:0] T358;
  wire[47:0] T359;
  wire[47:0] T360;
  wire[47:0] T361;
  wire[47:0] T362;
  wire[47:0] T363;
  wire[47:0] T364;
  wire[47:0] T365;
  wire[47:0] twiddle3_2_0_imag;
  wire[47:0] T366;
  wire[16:0] T367;
  wire[16:0] T368;
  wire[30:0] T369;
  wire T370;
  wire[47:0] T371;
  wire[47:0] T372;
  wire[47:0] T373;
  wire[46:0] twiddle3_2_1_imag;
  wire[46:0] T374;
  wire[42:0] T375;
  wire[42:0] T376;
  wire[3:0] T377;
  wire T378;
  wire[46:0] T379;
  wire[46:0] T380;
  wire T381;
  wire T382;
  wire[6:0] T383;
  wire[6:0] T384;
  wire[47:0] T385;
  wire[46:0] T386;
  wire[46:0] twiddle3_2_2_imag;
  wire[46:0] T387;
  wire[43:0] T388;
  wire[43:0] T389;
  wire[2:0] T390;
  wire T391;
  wire[46:0] T392;
  wire[46:0] T393;
  wire[46:0] twiddle3_2_3_imag;
  wire[46:0] T394;
  wire[44:0] T395;
  wire[44:0] T396;
  wire[1:0] T397;
  wire T398;
  wire[46:0] T399;
  wire[46:0] T400;
  wire T401;
  wire T402;
  wire T403;
  wire[47:0] T404;
  wire[46:0] T405;
  wire[46:0] T406;
  wire[46:0] twiddle3_2_4_imag;
  wire[46:0] T407;
  wire[44:0] T408;
  wire[44:0] T409;
  wire[1:0] T410;
  wire T411;
  wire[46:0] T412;
  wire[46:0] T413;
  wire[46:0] twiddle3_2_5_imag;
  wire[46:0] T414;
  wire[45:0] T415;
  wire[45:0] T416;
  wire T417;
  wire[46:0] T418;
  wire[46:0] T419;
  wire T420;
  wire[46:0] T421;
  wire[46:0] twiddle3_2_6_imag;
  wire[46:0] T422;
  wire[45:0] T423;
  wire[45:0] T424;
  wire T425;
  wire[46:0] T426;
  wire[46:0] T427;
  wire[46:0] twiddle3_2_7_imag;
  wire[46:0] T428;
  wire[45:0] T429;
  wire[45:0] T430;
  wire T431;
  wire[46:0] T432;
  wire[46:0] T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire[47:0] T438;
  wire[46:0] T439;
  wire[46:0] T440;
  wire[46:0] T441;
  wire[46:0] twiddle3_2_8_imag;
  wire[46:0] T442;
  wire[45:0] T443;
  wire[45:0] T444;
  wire T445;
  wire[46:0] T446;
  wire[46:0] T447;
  wire[46:0] twiddle3_2_9_imag;
  wire[46:0] T448;
  wire[45:0] T449;
  wire[45:0] T450;
  wire T451;
  wire[46:0] T452;
  wire[46:0] T453;
  wire T454;
  wire[46:0] T455;
  wire[46:0] twiddle3_2_10_imag;
  wire[46:0] T456;
  wire[45:0] T457;
  wire[45:0] T458;
  wire T459;
  wire[46:0] T460;
  wire[46:0] T461;
  wire[46:0] twiddle3_2_11_imag;
  wire[46:0] T462;
  wire[46:0] T463;
  wire[46:0] T464;
  wire[46:0] T465;
  wire T466;
  wire T467;
  wire[46:0] T468;
  wire[46:0] T469;
  wire[46:0] twiddle3_2_12_imag;
  wire[46:0] T470;
  wire[46:0] T471;
  wire[46:0] T472;
  wire[46:0] T473;
  wire[46:0] twiddle3_2_13_imag;
  wire[46:0] T474;
  wire[46:0] T475;
  wire[46:0] T476;
  wire[46:0] T477;
  wire T478;
  wire[46:0] T479;
  wire[46:0] twiddle3_2_14_imag;
  wire[46:0] T480;
  wire[46:0] T481;
  wire[46:0] T482;
  wire[46:0] T483;
  wire[46:0] twiddle3_2_15_imag;
  wire[46:0] T484;
  wire[46:0] T485;
  wire[46:0] T486;
  wire[46:0] T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire[47:0] T493;
  wire[46:0] T494;
  wire[46:0] T495;
  wire[46:0] T496;
  wire[46:0] T497;
  wire[46:0] twiddle3_2_16_imag;
  wire[46:0] T498;
  wire[46:0] T499;
  wire[46:0] T500;
  wire[46:0] T501;
  wire[46:0] twiddle3_2_17_imag;
  wire[46:0] T502;
  wire[46:0] T503;
  wire[46:0] T504;
  wire[46:0] T505;
  wire T506;
  wire[46:0] T507;
  wire[46:0] twiddle3_2_18_imag;
  wire[46:0] T508;
  wire[46:0] T509;
  wire[46:0] T510;
  wire[46:0] T511;
  wire[46:0] twiddle3_2_19_imag;
  wire[46:0] T512;
  wire[46:0] T513;
  wire[46:0] T514;
  wire[46:0] T515;
  wire T516;
  wire T517;
  wire[46:0] T518;
  wire[46:0] T519;
  wire[46:0] twiddle3_2_20_imag;
  wire[46:0] T520;
  wire[46:0] T521;
  wire[46:0] T522;
  wire[46:0] T523;
  wire[46:0] twiddle3_2_21_imag;
  wire[46:0] T524;
  wire[46:0] T525;
  wire[46:0] T526;
  wire[45:0] T527;
  wire[45:0] T528;
  wire T529;
  wire T530;
  wire[46:0] T531;
  wire[46:0] twiddle3_2_22_imag;
  wire[46:0] T532;
  wire[46:0] T533;
  wire[46:0] T534;
  wire[45:0] T535;
  wire[45:0] T536;
  wire T537;
  wire[46:0] twiddle3_2_23_imag;
  wire[46:0] T538;
  wire[46:0] T539;
  wire[46:0] T540;
  wire[45:0] T541;
  wire[45:0] T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire[46:0] T547;
  wire[46:0] T548;
  wire[46:0] T549;
  wire[46:0] twiddle3_2_24_imag;
  wire[46:0] T550;
  wire[46:0] T551;
  wire[46:0] T552;
  wire[45:0] T553;
  wire[45:0] T554;
  wire T555;
  wire[46:0] twiddle3_2_25_imag;
  wire[46:0] T556;
  wire[46:0] T557;
  wire[46:0] T558;
  wire[45:0] T559;
  wire[45:0] T560;
  wire T561;
  wire T562;
  wire[46:0] T563;
  wire[46:0] twiddle3_2_26_imag;
  wire[46:0] T564;
  wire[46:0] T565;
  wire[46:0] T566;
  wire[44:0] T567;
  wire[44:0] T568;
  wire[1:0] T569;
  wire T570;
  wire[46:0] twiddle3_2_27_imag;
  wire[46:0] T571;
  wire[46:0] T572;
  wire[46:0] T573;
  wire[44:0] T574;
  wire[44:0] T575;
  wire[1:0] T576;
  wire T577;
  wire T578;
  wire T579;
  wire[46:0] T580;
  wire[46:0] T581;
  wire[46:0] twiddle3_2_28_imag;
  wire[46:0] T582;
  wire[46:0] T583;
  wire[46:0] T584;
  wire[43:0] T585;
  wire[43:0] T586;
  wire[2:0] T587;
  wire T588;
  wire[46:0] twiddle3_2_29_imag;
  wire[46:0] T589;
  wire[46:0] T590;
  wire[46:0] T591;
  wire[43:0] T592;
  wire[43:0] T593;
  wire[2:0] T594;
  wire T595;
  wire T596;
  wire[46:0] T597;
  wire[46:0] twiddle3_2_30_imag;
  wire[46:0] T598;
  wire[46:0] T599;
  wire[46:0] T600;
  wire[41:0] T601;
  wire[41:0] T602;
  wire[4:0] T603;
  wire T604;
  wire[46:0] twiddle3_2_31_imag;
  wire[46:0] T605;
  wire[46:0] T606;
  wire[46:0] T607;
  wire[42:0] T608;
  wire[42:0] T609;
  wire[3:0] T610;
  wire T611;
  wire T612;
  wire T613;
  wire T614;
  wire T615;
  wire T616;
  wire T617;
  wire[47:0] T618;
  wire[46:0] T619;
  wire[46:0] T620;
  wire[46:0] T621;
  wire[46:0] T622;
  wire[46:0] T623;
  wire[46:0] twiddle3_2_32_imag;
  wire[46:0] T624;
  wire[46:0] T625;
  wire[46:0] T626;
  wire[43:0] T627;
  wire[43:0] T628;
  wire[2:0] T629;
  wire T630;
  wire[46:0] twiddle3_2_33_imag;
  wire[46:0] T631;
  wire[46:0] T632;
  wire[46:0] T633;
  wire[44:0] T634;
  wire[44:0] T635;
  wire[1:0] T636;
  wire T637;
  wire T638;
  wire[46:0] T639;
  wire[46:0] twiddle3_2_34_imag;
  wire[46:0] T640;
  wire[46:0] T641;
  wire[46:0] T642;
  wire[44:0] T643;
  wire[44:0] T644;
  wire[1:0] T645;
  wire T646;
  wire[46:0] twiddle3_2_35_imag;
  wire[46:0] T647;
  wire[46:0] T648;
  wire[46:0] T649;
  wire[44:0] T650;
  wire[44:0] T651;
  wire[1:0] T652;
  wire T653;
  wire T654;
  wire T655;
  wire[46:0] T656;
  wire[46:0] T657;
  wire[46:0] twiddle3_2_36_imag;
  wire[46:0] T658;
  wire[46:0] T659;
  wire[46:0] T660;
  wire[45:0] T661;
  wire[45:0] T662;
  wire T663;
  wire[46:0] twiddle3_2_37_imag;
  wire[46:0] T664;
  wire[46:0] T665;
  wire[46:0] T666;
  wire[45:0] T667;
  wire[45:0] T668;
  wire T669;
  wire T670;
  wire[46:0] T671;
  wire[46:0] twiddle3_2_38_imag;
  wire[46:0] T672;
  wire[46:0] T673;
  wire[46:0] T674;
  wire[45:0] T675;
  wire[45:0] T676;
  wire T677;
  wire[46:0] twiddle3_2_39_imag;
  wire[46:0] T678;
  wire[46:0] T679;
  wire[46:0] T680;
  wire[45:0] T681;
  wire[45:0] T682;
  wire T683;
  wire T684;
  wire T685;
  wire T686;
  wire[46:0] T687;
  wire[46:0] T688;
  wire[46:0] T689;
  wire[46:0] twiddle3_2_40_imag;
  wire[46:0] T690;
  wire[46:0] T691;
  wire[46:0] T692;
  wire[45:0] T693;
  wire[45:0] T694;
  wire T695;
  wire[46:0] twiddle3_2_41_imag;
  wire[46:0] T696;
  wire[46:0] T697;
  wire[46:0] T698;
  wire[46:0] T699;
  wire T700;
  wire[46:0] T701;
  wire[46:0] twiddle3_2_42_imag;
  wire[46:0] T702;
  wire[46:0] T703;
  wire[46:0] T704;
  wire[46:0] T705;
  wire[46:0] twiddle3_2_43_imag;
  wire[46:0] T706;
  wire[46:0] T707;
  wire[46:0] T708;
  wire[46:0] T709;
  wire T710;
  wire T711;
  wire[46:0] T712;
  wire[46:0] T713;
  wire[46:0] twiddle3_2_44_imag;
  wire[46:0] T714;
  wire[46:0] T715;
  wire[46:0] T716;
  wire[46:0] T717;
  wire[46:0] twiddle3_2_45_imag;
  wire[46:0] T718;
  wire[46:0] T719;
  wire[46:0] T720;
  wire[46:0] T721;
  wire T722;
  wire[46:0] T723;
  wire[46:0] twiddle3_2_46_imag;
  wire[46:0] T724;
  wire[46:0] T725;
  wire[46:0] T726;
  wire[46:0] T727;
  wire[46:0] twiddle3_2_47_imag;
  wire[46:0] T728;
  wire[46:0] T729;
  wire[46:0] T730;
  wire[46:0] T731;
  wire T732;
  wire T733;
  wire T734;
  wire T735;
  wire[46:0] T736;
  wire[46:0] T737;
  wire[46:0] T738;
  wire[46:0] T739;
  wire[46:0] twiddle3_2_48_imag;
  wire[46:0] T740;
  wire[46:0] T741;
  wire[46:0] T742;
  wire[46:0] T743;
  wire[46:0] twiddle3_2_49_imag;
  wire[46:0] T744;
  wire[46:0] T745;
  wire[46:0] T746;
  wire[46:0] T747;
  wire T748;
  wire[46:0] T749;
  wire[46:0] twiddle3_2_50_imag;
  wire[46:0] T750;
  wire[46:0] T751;
  wire[46:0] T752;
  wire[46:0] T753;
  wire[46:0] twiddle3_2_51_imag;
  wire[46:0] T754;
  wire[45:0] T755;
  wire[45:0] T756;
  wire T757;
  wire[46:0] T758;
  wire[46:0] T759;
  wire T760;
  wire T761;
  wire[46:0] T762;
  wire[46:0] T763;
  wire[46:0] twiddle3_2_52_imag;
  wire[46:0] T764;
  wire[45:0] T765;
  wire[45:0] T766;
  wire T767;
  wire[46:0] T768;
  wire[46:0] T769;
  wire[46:0] twiddle3_2_53_imag;
  wire[46:0] T770;
  wire[45:0] T771;
  wire[45:0] T772;
  wire T773;
  wire[46:0] T774;
  wire[46:0] T775;
  wire T776;
  wire[46:0] T777;
  wire[46:0] twiddle3_2_54_imag;
  wire[46:0] T778;
  wire[45:0] T779;
  wire[45:0] T780;
  wire T781;
  wire[46:0] T782;
  wire[46:0] T783;
  wire[46:0] twiddle3_2_55_imag;
  wire[46:0] T784;
  wire[45:0] T785;
  wire[45:0] T786;
  wire T787;
  wire[46:0] T788;
  wire[46:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire[46:0] T793;
  wire[46:0] T794;
  wire[46:0] T795;
  wire[46:0] twiddle3_2_56_imag;
  wire[46:0] T796;
  wire[44:0] T797;
  wire[44:0] T798;
  wire[1:0] T799;
  wire T800;
  wire[46:0] T801;
  wire[46:0] T802;
  wire[46:0] twiddle3_2_57_imag;
  wire[46:0] T803;
  wire[44:0] T804;
  wire[44:0] T805;
  wire[1:0] T806;
  wire T807;
  wire[46:0] T808;
  wire[46:0] T809;
  wire T810;
  wire[46:0] T811;
  wire[46:0] twiddle3_2_58_imag;
  wire[46:0] T812;
  wire[44:0] T813;
  wire[44:0] T814;
  wire[1:0] T815;
  wire T816;
  wire[46:0] T817;
  wire[46:0] T818;
  wire[46:0] twiddle3_2_59_imag;
  wire[46:0] T819;
  wire[43:0] T820;
  wire[43:0] T821;
  wire[2:0] T822;
  wire T823;
  wire[46:0] T824;
  wire[46:0] T825;
  wire T826;
  wire T827;
  wire[46:0] T828;
  wire[46:0] T829;
  wire[46:0] twiddle3_2_60_imag;
  wire[46:0] T830;
  wire[42:0] T831;
  wire[42:0] T832;
  wire[3:0] T833;
  wire T834;
  wire[46:0] T835;
  wire[46:0] T836;
  wire[46:0] twiddle3_2_61_imag;
  wire[46:0] T837;
  wire[40:0] T838;
  wire[40:0] T839;
  wire[5:0] T840;
  wire T841;
  wire[46:0] T842;
  wire[46:0] T843;
  wire T844;
  wire[46:0] T845;
  wire[46:0] twiddle3_2_62_imag;
  wire[46:0] T846;
  wire[43:0] T847;
  wire[43:0] T848;
  wire[2:0] T849;
  wire T850;
  wire[46:0] T851;
  wire[46:0] T852;
  wire[46:0] twiddle3_2_63_imag;
  wire[46:0] T853;
  wire[43:0] T854;
  wire[43:0] T855;
  wire[2:0] T856;
  wire T857;
  wire[46:0] T858;
  wire[46:0] T859;
  wire T860;
  wire T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire[47:0] T867;
  wire[46:0] T868;
  wire[46:0] T869;
  wire[46:0] T870;
  wire[46:0] T871;
  wire[46:0] T872;
  wire[46:0] twiddle3_2_64_imag;
  wire[46:0] T873;
  wire[44:0] T874;
  wire[44:0] T875;
  wire[1:0] T876;
  wire T877;
  wire[46:0] T878;
  wire[46:0] T879;
  wire[46:0] twiddle3_2_65_imag;
  wire[46:0] T880;
  wire[44:0] T881;
  wire[44:0] T882;
  wire[1:0] T883;
  wire T884;
  wire[46:0] T885;
  wire[46:0] T886;
  wire T887;
  wire[46:0] T888;
  wire[46:0] twiddle3_2_66_imag;
  wire[46:0] T889;
  wire[45:0] T890;
  wire[45:0] T891;
  wire T892;
  wire[46:0] T893;
  wire[46:0] T894;
  wire[46:0] twiddle3_2_67_imag;
  wire[46:0] T895;
  wire[45:0] T896;
  wire[45:0] T897;
  wire T898;
  wire[46:0] T899;
  wire[46:0] T900;
  wire T901;
  wire T902;
  wire[46:0] T903;
  wire[46:0] T904;
  wire[46:0] twiddle3_2_68_imag;
  wire[46:0] T905;
  wire[45:0] T906;
  wire[45:0] T907;
  wire T908;
  wire[46:0] T909;
  wire[46:0] T910;
  wire[46:0] twiddle3_2_69_imag;
  wire[46:0] T911;
  wire[45:0] T912;
  wire[45:0] T913;
  wire T914;
  wire[46:0] T915;
  wire[46:0] T916;
  wire T917;
  wire[46:0] T918;
  wire[46:0] twiddle3_2_70_imag;
  wire[46:0] T919;
  wire[45:0] T920;
  wire[45:0] T921;
  wire T922;
  wire[46:0] T923;
  wire[46:0] T924;
  wire[46:0] twiddle3_2_71_imag;
  wire[46:0] T925;
  wire[46:0] T926;
  wire[46:0] T927;
  wire[46:0] T928;
  wire T929;
  wire T930;
  wire T931;
  wire[46:0] T932;
  wire[46:0] T933;
  wire[46:0] T934;
  wire[46:0] twiddle3_2_72_imag;
  wire[46:0] T935;
  wire[46:0] T936;
  wire[46:0] T937;
  wire[46:0] T938;
  wire[46:0] twiddle3_2_73_imag;
  wire[46:0] T939;
  wire[46:0] T940;
  wire[46:0] T941;
  wire[46:0] T942;
  wire T943;
  wire[46:0] T944;
  wire[46:0] twiddle3_2_74_imag;
  wire[46:0] T945;
  wire[46:0] T946;
  wire[46:0] T947;
  wire[46:0] T948;
  wire[46:0] twiddle3_2_75_imag;
  wire[46:0] T949;
  wire[46:0] T950;
  wire[46:0] T951;
  wire[46:0] T952;
  wire T953;
  wire T954;
  wire[46:0] T955;
  wire[46:0] T956;
  wire[46:0] twiddle3_2_76_imag;
  wire[46:0] T957;
  wire[46:0] T958;
  wire[46:0] T959;
  wire[46:0] T960;
  wire[46:0] twiddle3_2_77_imag;
  wire[46:0] T961;
  wire[46:0] T962;
  wire[46:0] T963;
  wire[46:0] T964;
  wire T965;
  wire[46:0] T966;
  wire[46:0] twiddle3_2_78_imag;
  wire[46:0] T967;
  wire[46:0] T968;
  wire[46:0] T969;
  wire[46:0] T970;
  wire[46:0] twiddle3_2_79_imag;
  wire[46:0] T971;
  wire[46:0] T972;
  wire[46:0] T973;
  wire[46:0] T974;
  wire T975;
  wire T976;
  wire T977;
  wire T978;
  wire[46:0] twiddle3_2_80_imag;
  wire[46:0] T979;
  wire[46:0] T980;
  wire[46:0] T981;
  wire[46:0] T982;
  wire T983;
  wire T984;
  wire T985;
  wire[15:0] T986;
  wire[47:0] T987;
  wire[47:0] T988;
  wire[47:0] T989;
  wire[47:0] T990;
  wire[47:0] T991;
  wire[47:0] T992;
  wire[47:0] T993;
  wire[47:0] twiddle3_2_0_real;
  wire[47:0] T994;
  wire[16:0] T995;
  wire[16:0] T996;
  wire[30:0] T997;
  wire T998;
  wire[47:0] T999;
  wire[47:0] T1000;
  wire[47:0] T1001;
  wire[46:0] twiddle3_2_1_real;
  wire[46:0] T1002;
  wire[42:0] T1003;
  wire[42:0] T1004;
  wire[3:0] T1005;
  wire T1006;
  wire[46:0] T1007;
  wire[46:0] T1008;
  wire T1009;
  wire T1010;
  wire[47:0] T1011;
  wire[46:0] T1012;
  wire[46:0] twiddle3_2_2_real;
  wire[46:0] T1013;
  wire[43:0] T1014;
  wire[43:0] T1015;
  wire[2:0] T1016;
  wire T1017;
  wire[46:0] T1018;
  wire[46:0] T1019;
  wire[46:0] twiddle3_2_3_real;
  wire[46:0] T1020;
  wire[44:0] T1021;
  wire[44:0] T1022;
  wire[1:0] T1023;
  wire T1024;
  wire[46:0] T1025;
  wire[46:0] T1026;
  wire T1027;
  wire T1028;
  wire T1029;
  wire[47:0] T1030;
  wire[46:0] T1031;
  wire[46:0] T1032;
  wire[46:0] twiddle3_2_4_real;
  wire[46:0] T1033;
  wire[44:0] T1034;
  wire[44:0] T1035;
  wire[1:0] T1036;
  wire T1037;
  wire[46:0] T1038;
  wire[46:0] T1039;
  wire[46:0] twiddle3_2_5_real;
  wire[46:0] T1040;
  wire[45:0] T1041;
  wire[45:0] T1042;
  wire T1043;
  wire[46:0] T1044;
  wire[46:0] T1045;
  wire T1046;
  wire[46:0] T1047;
  wire[46:0] twiddle3_2_6_real;
  wire[46:0] T1048;
  wire[45:0] T1049;
  wire[45:0] T1050;
  wire T1051;
  wire[46:0] T1052;
  wire[46:0] T1053;
  wire[46:0] twiddle3_2_7_real;
  wire[46:0] T1054;
  wire[45:0] T1055;
  wire[45:0] T1056;
  wire T1057;
  wire[46:0] T1058;
  wire[46:0] T1059;
  wire T1060;
  wire T1061;
  wire T1062;
  wire T1063;
  wire[47:0] T1064;
  wire[46:0] T1065;
  wire[46:0] T1066;
  wire[46:0] T1067;
  wire[46:0] twiddle3_2_8_real;
  wire[46:0] T1068;
  wire[45:0] T1069;
  wire[45:0] T1070;
  wire T1071;
  wire[46:0] T1072;
  wire[46:0] T1073;
  wire[46:0] twiddle3_2_9_real;
  wire[46:0] T1074;
  wire[45:0] T1075;
  wire[45:0] T1076;
  wire T1077;
  wire[46:0] T1078;
  wire[46:0] T1079;
  wire T1080;
  wire[46:0] T1081;
  wire[46:0] twiddle3_2_10_real;
  wire[46:0] T1082;
  wire[45:0] T1083;
  wire[45:0] T1084;
  wire T1085;
  wire[46:0] T1086;
  wire[46:0] T1087;
  wire[46:0] twiddle3_2_11_real;
  wire[46:0] T1088;
  wire[46:0] T1089;
  wire[46:0] T1090;
  wire[46:0] T1091;
  wire T1092;
  wire T1093;
  wire[46:0] T1094;
  wire[46:0] T1095;
  wire[46:0] twiddle3_2_12_real;
  wire[46:0] T1096;
  wire[46:0] T1097;
  wire[46:0] T1098;
  wire[46:0] T1099;
  wire[46:0] twiddle3_2_13_real;
  wire[46:0] T1100;
  wire[46:0] T1101;
  wire[46:0] T1102;
  wire[46:0] T1103;
  wire T1104;
  wire[46:0] T1105;
  wire[46:0] twiddle3_2_14_real;
  wire[46:0] T1106;
  wire[46:0] T1107;
  wire[46:0] T1108;
  wire[46:0] T1109;
  wire[46:0] twiddle3_2_15_real;
  wire[46:0] T1110;
  wire[46:0] T1111;
  wire[46:0] T1112;
  wire[46:0] T1113;
  wire T1114;
  wire T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire[47:0] T1119;
  wire[46:0] T1120;
  wire[46:0] T1121;
  wire[46:0] T1122;
  wire[46:0] T1123;
  wire[46:0] twiddle3_2_16_real;
  wire[46:0] T1124;
  wire[46:0] T1125;
  wire[46:0] T1126;
  wire[46:0] T1127;
  wire[46:0] twiddle3_2_17_real;
  wire[46:0] T1128;
  wire[46:0] T1129;
  wire[46:0] T1130;
  wire[46:0] T1131;
  wire T1132;
  wire[46:0] T1133;
  wire[46:0] twiddle3_2_18_real;
  wire[46:0] T1134;
  wire[46:0] T1135;
  wire[46:0] T1136;
  wire[46:0] T1137;
  wire[46:0] twiddle3_2_19_real;
  wire[46:0] T1138;
  wire[46:0] T1139;
  wire[46:0] T1140;
  wire[46:0] T1141;
  wire T1142;
  wire T1143;
  wire[46:0] T1144;
  wire[46:0] T1145;
  wire[46:0] twiddle3_2_20_real;
  wire[46:0] T1146;
  wire[46:0] T1147;
  wire[46:0] T1148;
  wire[46:0] T1149;
  wire[46:0] twiddle3_2_21_real;
  wire[46:0] T1150;
  wire[46:0] T1151;
  wire[46:0] T1152;
  wire[45:0] T1153;
  wire[45:0] T1154;
  wire T1155;
  wire T1156;
  wire[46:0] T1157;
  wire[46:0] twiddle3_2_22_real;
  wire[46:0] T1158;
  wire[46:0] T1159;
  wire[46:0] T1160;
  wire[45:0] T1161;
  wire[45:0] T1162;
  wire T1163;
  wire[46:0] twiddle3_2_23_real;
  wire[46:0] T1164;
  wire[46:0] T1165;
  wire[46:0] T1166;
  wire[45:0] T1167;
  wire[45:0] T1168;
  wire T1169;
  wire T1170;
  wire T1171;
  wire T1172;
  wire[46:0] T1173;
  wire[46:0] T1174;
  wire[46:0] T1175;
  wire[46:0] twiddle3_2_24_real;
  wire[46:0] T1176;
  wire[46:0] T1177;
  wire[46:0] T1178;
  wire[45:0] T1179;
  wire[45:0] T1180;
  wire T1181;
  wire[46:0] twiddle3_2_25_real;
  wire[46:0] T1182;
  wire[46:0] T1183;
  wire[46:0] T1184;
  wire[45:0] T1185;
  wire[45:0] T1186;
  wire T1187;
  wire T1188;
  wire[46:0] T1189;
  wire[46:0] twiddle3_2_26_real;
  wire[46:0] T1190;
  wire[46:0] T1191;
  wire[46:0] T1192;
  wire[44:0] T1193;
  wire[44:0] T1194;
  wire[1:0] T1195;
  wire T1196;
  wire[46:0] twiddle3_2_27_real;
  wire[46:0] T1197;
  wire[46:0] T1198;
  wire[46:0] T1199;
  wire[44:0] T1200;
  wire[44:0] T1201;
  wire[1:0] T1202;
  wire T1203;
  wire T1204;
  wire T1205;
  wire[46:0] T1206;
  wire[46:0] T1207;
  wire[46:0] twiddle3_2_28_real;
  wire[46:0] T1208;
  wire[46:0] T1209;
  wire[46:0] T1210;
  wire[43:0] T1211;
  wire[43:0] T1212;
  wire[2:0] T1213;
  wire T1214;
  wire[46:0] twiddle3_2_29_real;
  wire[46:0] T1215;
  wire[46:0] T1216;
  wire[46:0] T1217;
  wire[43:0] T1218;
  wire[43:0] T1219;
  wire[2:0] T1220;
  wire T1221;
  wire T1222;
  wire[46:0] T1223;
  wire[46:0] twiddle3_2_30_real;
  wire[46:0] T1224;
  wire[46:0] T1225;
  wire[46:0] T1226;
  wire[41:0] T1227;
  wire[41:0] T1228;
  wire[4:0] T1229;
  wire T1230;
  wire[46:0] twiddle3_2_31_real;
  wire[46:0] T1231;
  wire[46:0] T1232;
  wire[46:0] T1233;
  wire[42:0] T1234;
  wire[42:0] T1235;
  wire[3:0] T1236;
  wire T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire[47:0] T1244;
  wire[46:0] T1245;
  wire[46:0] T1246;
  wire[46:0] T1247;
  wire[46:0] T1248;
  wire[46:0] T1249;
  wire[46:0] twiddle3_2_32_real;
  wire[46:0] T1250;
  wire[46:0] T1251;
  wire[46:0] T1252;
  wire[43:0] T1253;
  wire[43:0] T1254;
  wire[2:0] T1255;
  wire T1256;
  wire[46:0] twiddle3_2_33_real;
  wire[46:0] T1257;
  wire[46:0] T1258;
  wire[46:0] T1259;
  wire[44:0] T1260;
  wire[44:0] T1261;
  wire[1:0] T1262;
  wire T1263;
  wire T1264;
  wire[46:0] T1265;
  wire[46:0] twiddle3_2_34_real;
  wire[46:0] T1266;
  wire[46:0] T1267;
  wire[46:0] T1268;
  wire[44:0] T1269;
  wire[44:0] T1270;
  wire[1:0] T1271;
  wire T1272;
  wire[46:0] twiddle3_2_35_real;
  wire[46:0] T1273;
  wire[46:0] T1274;
  wire[46:0] T1275;
  wire[44:0] T1276;
  wire[44:0] T1277;
  wire[1:0] T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  wire[46:0] T1282;
  wire[46:0] T1283;
  wire[46:0] twiddle3_2_36_real;
  wire[46:0] T1284;
  wire[46:0] T1285;
  wire[46:0] T1286;
  wire[45:0] T1287;
  wire[45:0] T1288;
  wire T1289;
  wire[46:0] twiddle3_2_37_real;
  wire[46:0] T1290;
  wire[46:0] T1291;
  wire[46:0] T1292;
  wire[45:0] T1293;
  wire[45:0] T1294;
  wire T1295;
  wire T1296;
  wire[46:0] T1297;
  wire[46:0] twiddle3_2_38_real;
  wire[46:0] T1298;
  wire[46:0] T1299;
  wire[46:0] T1300;
  wire[45:0] T1301;
  wire[45:0] T1302;
  wire T1303;
  wire[46:0] twiddle3_2_39_real;
  wire[46:0] T1304;
  wire[46:0] T1305;
  wire[46:0] T1306;
  wire[45:0] T1307;
  wire[45:0] T1308;
  wire T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire[46:0] T1313;
  wire[46:0] T1314;
  wire[46:0] T1315;
  wire[46:0] twiddle3_2_40_real;
  wire[46:0] T1316;
  wire[46:0] T1317;
  wire[46:0] T1318;
  wire[45:0] T1319;
  wire[45:0] T1320;
  wire T1321;
  wire[46:0] twiddle3_2_41_real;
  wire[46:0] T1322;
  wire[46:0] T1323;
  wire[46:0] T1324;
  wire[46:0] T1325;
  wire T1326;
  wire[46:0] T1327;
  wire[46:0] twiddle3_2_42_real;
  wire[46:0] T1328;
  wire[46:0] T1329;
  wire[46:0] T1330;
  wire[46:0] T1331;
  wire[46:0] twiddle3_2_43_real;
  wire[46:0] T1332;
  wire[46:0] T1333;
  wire[46:0] T1334;
  wire[46:0] T1335;
  wire T1336;
  wire T1337;
  wire[46:0] T1338;
  wire[46:0] T1339;
  wire[46:0] twiddle3_2_44_real;
  wire[46:0] T1340;
  wire[46:0] T1341;
  wire[46:0] T1342;
  wire[46:0] T1343;
  wire[46:0] twiddle3_2_45_real;
  wire[46:0] T1344;
  wire[46:0] T1345;
  wire[46:0] T1346;
  wire[46:0] T1347;
  wire T1348;
  wire[46:0] T1349;
  wire[46:0] twiddle3_2_46_real;
  wire[46:0] T1350;
  wire[46:0] T1351;
  wire[46:0] T1352;
  wire[46:0] T1353;
  wire[46:0] twiddle3_2_47_real;
  wire[46:0] T1354;
  wire[46:0] T1355;
  wire[46:0] T1356;
  wire[46:0] T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire T1361;
  wire[46:0] T1362;
  wire[46:0] T1363;
  wire[46:0] T1364;
  wire[46:0] T1365;
  wire[46:0] twiddle3_2_48_real;
  wire[46:0] T1366;
  wire[46:0] T1367;
  wire[46:0] T1368;
  wire[46:0] T1369;
  wire[46:0] twiddle3_2_49_real;
  wire[46:0] T1370;
  wire[46:0] T1371;
  wire[46:0] T1372;
  wire[46:0] T1373;
  wire T1374;
  wire[46:0] T1375;
  wire[46:0] twiddle3_2_50_real;
  wire[46:0] T1376;
  wire[46:0] T1377;
  wire[46:0] T1378;
  wire[46:0] T1379;
  wire[46:0] twiddle3_2_51_real;
  wire[46:0] T1380;
  wire[45:0] T1381;
  wire[45:0] T1382;
  wire T1383;
  wire[46:0] T1384;
  wire[46:0] T1385;
  wire T1386;
  wire T1387;
  wire[46:0] T1388;
  wire[46:0] T1389;
  wire[46:0] twiddle3_2_52_real;
  wire[46:0] T1390;
  wire[45:0] T1391;
  wire[45:0] T1392;
  wire T1393;
  wire[46:0] T1394;
  wire[46:0] T1395;
  wire[46:0] twiddle3_2_53_real;
  wire[46:0] T1396;
  wire[45:0] T1397;
  wire[45:0] T1398;
  wire T1399;
  wire[46:0] T1400;
  wire[46:0] T1401;
  wire T1402;
  wire[46:0] T1403;
  wire[46:0] twiddle3_2_54_real;
  wire[46:0] T1404;
  wire[45:0] T1405;
  wire[45:0] T1406;
  wire T1407;
  wire[46:0] T1408;
  wire[46:0] T1409;
  wire[46:0] twiddle3_2_55_real;
  wire[46:0] T1410;
  wire[45:0] T1411;
  wire[45:0] T1412;
  wire T1413;
  wire[46:0] T1414;
  wire[46:0] T1415;
  wire T1416;
  wire T1417;
  wire T1418;
  wire[46:0] T1419;
  wire[46:0] T1420;
  wire[46:0] T1421;
  wire[46:0] twiddle3_2_56_real;
  wire[46:0] T1422;
  wire[44:0] T1423;
  wire[44:0] T1424;
  wire[1:0] T1425;
  wire T1426;
  wire[46:0] T1427;
  wire[46:0] T1428;
  wire[46:0] twiddle3_2_57_real;
  wire[46:0] T1429;
  wire[44:0] T1430;
  wire[44:0] T1431;
  wire[1:0] T1432;
  wire T1433;
  wire[46:0] T1434;
  wire[46:0] T1435;
  wire T1436;
  wire[46:0] T1437;
  wire[46:0] twiddle3_2_58_real;
  wire[46:0] T1438;
  wire[44:0] T1439;
  wire[44:0] T1440;
  wire[1:0] T1441;
  wire T1442;
  wire[46:0] T1443;
  wire[46:0] T1444;
  wire[46:0] twiddle3_2_59_real;
  wire[46:0] T1445;
  wire[43:0] T1446;
  wire[43:0] T1447;
  wire[2:0] T1448;
  wire T1449;
  wire[46:0] T1450;
  wire[46:0] T1451;
  wire T1452;
  wire T1453;
  wire[46:0] T1454;
  wire[46:0] T1455;
  wire[46:0] twiddle3_2_60_real;
  wire[46:0] T1456;
  wire[42:0] T1457;
  wire[42:0] T1458;
  wire[3:0] T1459;
  wire T1460;
  wire[46:0] T1461;
  wire[46:0] T1462;
  wire[46:0] twiddle3_2_61_real;
  wire[46:0] T1463;
  wire[40:0] T1464;
  wire[40:0] T1465;
  wire[5:0] T1466;
  wire T1467;
  wire[46:0] T1468;
  wire[46:0] T1469;
  wire T1470;
  wire[46:0] T1471;
  wire[46:0] twiddle3_2_62_real;
  wire[46:0] T1472;
  wire[43:0] T1473;
  wire[43:0] T1474;
  wire[2:0] T1475;
  wire T1476;
  wire[46:0] T1477;
  wire[46:0] T1478;
  wire[46:0] twiddle3_2_63_real;
  wire[46:0] T1479;
  wire[43:0] T1480;
  wire[43:0] T1481;
  wire[2:0] T1482;
  wire T1483;
  wire[46:0] T1484;
  wire[46:0] T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire T1489;
  wire T1490;
  wire T1491;
  wire T1492;
  wire[47:0] T1493;
  wire[46:0] T1494;
  wire[46:0] T1495;
  wire[46:0] T1496;
  wire[46:0] T1497;
  wire[46:0] T1498;
  wire[46:0] twiddle3_2_64_real;
  wire[46:0] T1499;
  wire[44:0] T1500;
  wire[44:0] T1501;
  wire[1:0] T1502;
  wire T1503;
  wire[46:0] T1504;
  wire[46:0] T1505;
  wire[46:0] twiddle3_2_65_real;
  wire[46:0] T1506;
  wire[44:0] T1507;
  wire[44:0] T1508;
  wire[1:0] T1509;
  wire T1510;
  wire[46:0] T1511;
  wire[46:0] T1512;
  wire T1513;
  wire[46:0] T1514;
  wire[46:0] twiddle3_2_66_real;
  wire[46:0] T1515;
  wire[45:0] T1516;
  wire[45:0] T1517;
  wire T1518;
  wire[46:0] T1519;
  wire[46:0] T1520;
  wire[46:0] twiddle3_2_67_real;
  wire[46:0] T1521;
  wire[45:0] T1522;
  wire[45:0] T1523;
  wire T1524;
  wire[46:0] T1525;
  wire[46:0] T1526;
  wire T1527;
  wire T1528;
  wire[46:0] T1529;
  wire[46:0] T1530;
  wire[46:0] twiddle3_2_68_real;
  wire[46:0] T1531;
  wire[45:0] T1532;
  wire[45:0] T1533;
  wire T1534;
  wire[46:0] T1535;
  wire[46:0] T1536;
  wire[46:0] twiddle3_2_69_real;
  wire[46:0] T1537;
  wire[45:0] T1538;
  wire[45:0] T1539;
  wire T1540;
  wire[46:0] T1541;
  wire[46:0] T1542;
  wire T1543;
  wire[46:0] T1544;
  wire[46:0] twiddle3_2_70_real;
  wire[46:0] T1545;
  wire[45:0] T1546;
  wire[45:0] T1547;
  wire T1548;
  wire[46:0] T1549;
  wire[46:0] T1550;
  wire[46:0] twiddle3_2_71_real;
  wire[46:0] T1551;
  wire[46:0] T1552;
  wire[46:0] T1553;
  wire[46:0] T1554;
  wire T1555;
  wire T1556;
  wire T1557;
  wire[46:0] T1558;
  wire[46:0] T1559;
  wire[46:0] T1560;
  wire[46:0] twiddle3_2_72_real;
  wire[46:0] T1561;
  wire[46:0] T1562;
  wire[46:0] T1563;
  wire[46:0] T1564;
  wire[46:0] twiddle3_2_73_real;
  wire[46:0] T1565;
  wire[46:0] T1566;
  wire[46:0] T1567;
  wire[46:0] T1568;
  wire T1569;
  wire[46:0] T1570;
  wire[46:0] twiddle3_2_74_real;
  wire[46:0] T1571;
  wire[46:0] T1572;
  wire[46:0] T1573;
  wire[46:0] T1574;
  wire[46:0] twiddle3_2_75_real;
  wire[46:0] T1575;
  wire[46:0] T1576;
  wire[46:0] T1577;
  wire[46:0] T1578;
  wire T1579;
  wire T1580;
  wire[46:0] T1581;
  wire[46:0] T1582;
  wire[46:0] twiddle3_2_76_real;
  wire[46:0] T1583;
  wire[46:0] T1584;
  wire[46:0] T1585;
  wire[46:0] T1586;
  wire[46:0] twiddle3_2_77_real;
  wire[46:0] T1587;
  wire[46:0] T1588;
  wire[46:0] T1589;
  wire[46:0] T1590;
  wire T1591;
  wire[46:0] T1592;
  wire[46:0] twiddle3_2_78_real;
  wire[46:0] T1593;
  wire[46:0] T1594;
  wire[46:0] T1595;
  wire[46:0] T1596;
  wire[46:0] twiddle3_2_79_real;
  wire[46:0] T1597;
  wire[46:0] T1598;
  wire[46:0] T1599;
  wire[46:0] T1600;
  wire T1601;
  wire T1602;
  wire T1603;
  wire T1604;
  wire[46:0] twiddle3_2_80_real;
  wire[46:0] T1605;
  wire[46:0] T1606;
  wire[46:0] T1607;
  wire[46:0] T1608;
  wire T1609;
  wire T1610;
  wire T1611;
  wire[15:0] T1612;
  wire[47:0] T1613;
  wire[47:0] T1614;
  wire[47:0] T1615;
  wire[47:0] T1616;
  wire[47:0] T1617;
  wire[47:0] T1618;
  wire[47:0] T1619;
  wire[47:0] twiddle3_1_0_imag;
  wire[47:0] T1620;
  wire[16:0] T1621;
  wire[16:0] T1622;
  wire[30:0] T1623;
  wire T1624;
  wire[47:0] T1625;
  wire[47:0] T1626;
  wire[47:0] T1627;
  wire[46:0] twiddle3_1_1_imag;
  wire[46:0] T1628;
  wire[41:0] T1629;
  wire[41:0] T1630;
  wire[4:0] T1631;
  wire T1632;
  wire[46:0] T1633;
  wire[46:0] T1634;
  wire T1635;
  wire T1636;
  wire[6:0] T1637;
  wire[6:0] T1638;
  wire[47:0] T1639;
  wire[46:0] T1640;
  wire[46:0] twiddle3_1_2_imag;
  wire[46:0] T1641;
  wire[42:0] T1642;
  wire[42:0] T1643;
  wire[3:0] T1644;
  wire T1645;
  wire[46:0] T1646;
  wire[46:0] T1647;
  wire[46:0] twiddle3_1_3_imag;
  wire[46:0] T1648;
  wire[43:0] T1649;
  wire[43:0] T1650;
  wire[2:0] T1651;
  wire T1652;
  wire[46:0] T1653;
  wire[46:0] T1654;
  wire T1655;
  wire T1656;
  wire T1657;
  wire[47:0] T1658;
  wire[46:0] T1659;
  wire[46:0] T1660;
  wire[46:0] twiddle3_1_4_imag;
  wire[46:0] T1661;
  wire[43:0] T1662;
  wire[43:0] T1663;
  wire[2:0] T1664;
  wire T1665;
  wire[46:0] T1666;
  wire[46:0] T1667;
  wire[46:0] twiddle3_1_5_imag;
  wire[46:0] T1668;
  wire[44:0] T1669;
  wire[44:0] T1670;
  wire[1:0] T1671;
  wire T1672;
  wire[46:0] T1673;
  wire[46:0] T1674;
  wire T1675;
  wire[46:0] T1676;
  wire[46:0] twiddle3_1_6_imag;
  wire[46:0] T1677;
  wire[44:0] T1678;
  wire[44:0] T1679;
  wire[1:0] T1680;
  wire T1681;
  wire[46:0] T1682;
  wire[46:0] T1683;
  wire[46:0] twiddle3_1_7_imag;
  wire[46:0] T1684;
  wire[44:0] T1685;
  wire[44:0] T1686;
  wire[1:0] T1687;
  wire T1688;
  wire[46:0] T1689;
  wire[46:0] T1690;
  wire T1691;
  wire T1692;
  wire T1693;
  wire T1694;
  wire[47:0] T1695;
  wire[46:0] T1696;
  wire[46:0] T1697;
  wire[46:0] T1698;
  wire[46:0] twiddle3_1_8_imag;
  wire[46:0] T1699;
  wire[44:0] T1700;
  wire[44:0] T1701;
  wire[1:0] T1702;
  wire T1703;
  wire[46:0] T1704;
  wire[46:0] T1705;
  wire[46:0] twiddle3_1_9_imag;
  wire[46:0] T1706;
  wire[44:0] T1707;
  wire[44:0] T1708;
  wire[1:0] T1709;
  wire T1710;
  wire[46:0] T1711;
  wire[46:0] T1712;
  wire T1713;
  wire[46:0] T1714;
  wire[46:0] twiddle3_1_10_imag;
  wire[46:0] T1715;
  wire[45:0] T1716;
  wire[45:0] T1717;
  wire T1718;
  wire[46:0] T1719;
  wire[46:0] T1720;
  wire[46:0] twiddle3_1_11_imag;
  wire[46:0] T1721;
  wire[45:0] T1722;
  wire[45:0] T1723;
  wire T1724;
  wire[46:0] T1725;
  wire[46:0] T1726;
  wire T1727;
  wire T1728;
  wire[46:0] T1729;
  wire[46:0] T1730;
  wire[46:0] twiddle3_1_12_imag;
  wire[46:0] T1731;
  wire[45:0] T1732;
  wire[45:0] T1733;
  wire T1734;
  wire[46:0] T1735;
  wire[46:0] T1736;
  wire[46:0] twiddle3_1_13_imag;
  wire[46:0] T1737;
  wire[45:0] T1738;
  wire[45:0] T1739;
  wire T1740;
  wire[46:0] T1741;
  wire[46:0] T1742;
  wire T1743;
  wire[46:0] T1744;
  wire[46:0] twiddle3_1_14_imag;
  wire[46:0] T1745;
  wire[45:0] T1746;
  wire[45:0] T1747;
  wire T1748;
  wire[46:0] T1749;
  wire[46:0] T1750;
  wire[46:0] twiddle3_1_15_imag;
  wire[46:0] T1751;
  wire[45:0] T1752;
  wire[45:0] T1753;
  wire T1754;
  wire[46:0] T1755;
  wire[46:0] T1756;
  wire T1757;
  wire T1758;
  wire T1759;
  wire T1760;
  wire T1761;
  wire[47:0] T1762;
  wire[46:0] T1763;
  wire[46:0] T1764;
  wire[46:0] T1765;
  wire[46:0] T1766;
  wire[46:0] twiddle3_1_16_imag;
  wire[46:0] T1767;
  wire[45:0] T1768;
  wire[45:0] T1769;
  wire T1770;
  wire[46:0] T1771;
  wire[46:0] T1772;
  wire[46:0] twiddle3_1_17_imag;
  wire[46:0] T1773;
  wire[45:0] T1774;
  wire[45:0] T1775;
  wire T1776;
  wire[46:0] T1777;
  wire[46:0] T1778;
  wire T1779;
  wire[46:0] T1780;
  wire[46:0] twiddle3_1_18_imag;
  wire[46:0] T1781;
  wire[45:0] T1782;
  wire[45:0] T1783;
  wire T1784;
  wire[46:0] T1785;
  wire[46:0] T1786;
  wire[46:0] twiddle3_1_19_imag;
  wire[46:0] T1787;
  wire[45:0] T1788;
  wire[45:0] T1789;
  wire T1790;
  wire[46:0] T1791;
  wire[46:0] T1792;
  wire T1793;
  wire T1794;
  wire[46:0] T1795;
  wire[46:0] T1796;
  wire[46:0] twiddle3_1_20_imag;
  wire[46:0] T1797;
  wire[45:0] T1798;
  wire[45:0] T1799;
  wire T1800;
  wire[46:0] T1801;
  wire[46:0] T1802;
  wire[46:0] twiddle3_1_21_imag;
  wire[46:0] T1803;
  wire[46:0] T1804;
  wire[46:0] T1805;
  wire[46:0] T1806;
  wire T1807;
  wire[46:0] T1808;
  wire[46:0] twiddle3_1_22_imag;
  wire[46:0] T1809;
  wire[46:0] T1810;
  wire[46:0] T1811;
  wire[46:0] T1812;
  wire[46:0] twiddle3_1_23_imag;
  wire[46:0] T1813;
  wire[46:0] T1814;
  wire[46:0] T1815;
  wire[46:0] T1816;
  wire T1817;
  wire T1818;
  wire T1819;
  wire[46:0] T1820;
  wire[46:0] T1821;
  wire[46:0] T1822;
  wire[46:0] twiddle3_1_24_imag;
  wire[46:0] T1823;
  wire[46:0] T1824;
  wire[46:0] T1825;
  wire[46:0] T1826;
  wire[46:0] twiddle3_1_25_imag;
  wire[46:0] T1827;
  wire[46:0] T1828;
  wire[46:0] T1829;
  wire[46:0] T1830;
  wire T1831;
  wire[46:0] T1832;
  wire[46:0] twiddle3_1_26_imag;
  wire[46:0] T1833;
  wire[46:0] T1834;
  wire[46:0] T1835;
  wire[46:0] T1836;
  wire[46:0] twiddle3_1_27_imag;
  wire[46:0] T1837;
  wire[46:0] T1838;
  wire[46:0] T1839;
  wire[46:0] T1840;
  wire T1841;
  wire T1842;
  wire[46:0] T1843;
  wire[46:0] T1844;
  wire[46:0] twiddle3_1_28_imag;
  wire[46:0] T1845;
  wire[46:0] T1846;
  wire[46:0] T1847;
  wire[46:0] T1848;
  wire[46:0] twiddle3_1_29_imag;
  wire[46:0] T1849;
  wire[46:0] T1850;
  wire[46:0] T1851;
  wire[46:0] T1852;
  wire T1853;
  wire[46:0] T1854;
  wire[46:0] twiddle3_1_30_imag;
  wire[46:0] T1855;
  wire[46:0] T1856;
  wire[46:0] T1857;
  wire[46:0] T1858;
  wire[46:0] twiddle3_1_31_imag;
  wire[46:0] T1859;
  wire[46:0] T1860;
  wire[46:0] T1861;
  wire[46:0] T1862;
  wire T1863;
  wire T1864;
  wire T1865;
  wire T1866;
  wire T1867;
  wire T1868;
  wire[47:0] T1869;
  wire[46:0] T1870;
  wire[46:0] T1871;
  wire[46:0] T1872;
  wire[46:0] T1873;
  wire[46:0] T1874;
  wire[46:0] twiddle3_1_32_imag;
  wire[46:0] T1875;
  wire[46:0] T1876;
  wire[46:0] T1877;
  wire[46:0] T1878;
  wire[46:0] twiddle3_1_33_imag;
  wire[46:0] T1879;
  wire[46:0] T1880;
  wire[46:0] T1881;
  wire[46:0] T1882;
  wire T1883;
  wire[46:0] T1884;
  wire[46:0] twiddle3_1_34_imag;
  wire[46:0] T1885;
  wire[46:0] T1886;
  wire[46:0] T1887;
  wire[46:0] T1888;
  wire[46:0] twiddle3_1_35_imag;
  wire[46:0] T1889;
  wire[46:0] T1890;
  wire[46:0] T1891;
  wire[46:0] T1892;
  wire T1893;
  wire T1894;
  wire[46:0] T1895;
  wire[46:0] T1896;
  wire[46:0] twiddle3_1_36_imag;
  wire[46:0] T1897;
  wire[46:0] T1898;
  wire[46:0] T1899;
  wire[46:0] T1900;
  wire[46:0] twiddle3_1_37_imag;
  wire[46:0] T1901;
  wire[46:0] T1902;
  wire[46:0] T1903;
  wire[46:0] T1904;
  wire T1905;
  wire[46:0] T1906;
  wire[46:0] twiddle3_1_38_imag;
  wire[46:0] T1907;
  wire[46:0] T1908;
  wire[46:0] T1909;
  wire[46:0] T1910;
  wire[46:0] twiddle3_1_39_imag;
  wire[46:0] T1911;
  wire[46:0] T1912;
  wire[46:0] T1913;
  wire[46:0] T1914;
  wire T1915;
  wire T1916;
  wire T1917;
  wire[46:0] T1918;
  wire[46:0] T1919;
  wire[46:0] T1920;
  wire[46:0] twiddle3_1_40_imag;
  wire[46:0] T1921;
  wire[46:0] T1922;
  wire[46:0] T1923;
  wire[46:0] T1924;
  wire[46:0] twiddle3_1_41_imag;
  wire[46:0] T1925;
  wire[46:0] T1926;
  wire[46:0] T1927;
  wire[45:0] T1928;
  wire[45:0] T1929;
  wire T1930;
  wire T1931;
  wire[46:0] T1932;
  wire[46:0] twiddle3_1_42_imag;
  wire[46:0] T1933;
  wire[46:0] T1934;
  wire[46:0] T1935;
  wire[45:0] T1936;
  wire[45:0] T1937;
  wire T1938;
  wire[46:0] twiddle3_1_43_imag;
  wire[46:0] T1939;
  wire[46:0] T1940;
  wire[46:0] T1941;
  wire[45:0] T1942;
  wire[45:0] T1943;
  wire T1944;
  wire T1945;
  wire T1946;
  wire[46:0] T1947;
  wire[46:0] T1948;
  wire[46:0] twiddle3_1_44_imag;
  wire[46:0] T1949;
  wire[46:0] T1950;
  wire[46:0] T1951;
  wire[45:0] T1952;
  wire[45:0] T1953;
  wire T1954;
  wire[46:0] twiddle3_1_45_imag;
  wire[46:0] T1955;
  wire[46:0] T1956;
  wire[46:0] T1957;
  wire[45:0] T1958;
  wire[45:0] T1959;
  wire T1960;
  wire T1961;
  wire[46:0] T1962;
  wire[46:0] twiddle3_1_46_imag;
  wire[46:0] T1963;
  wire[46:0] T1964;
  wire[46:0] T1965;
  wire[45:0] T1966;
  wire[45:0] T1967;
  wire T1968;
  wire[46:0] twiddle3_1_47_imag;
  wire[46:0] T1969;
  wire[46:0] T1970;
  wire[46:0] T1971;
  wire[45:0] T1972;
  wire[45:0] T1973;
  wire T1974;
  wire T1975;
  wire T1976;
  wire T1977;
  wire T1978;
  wire[46:0] T1979;
  wire[46:0] T1980;
  wire[46:0] T1981;
  wire[46:0] T1982;
  wire[46:0] twiddle3_1_48_imag;
  wire[46:0] T1983;
  wire[46:0] T1984;
  wire[46:0] T1985;
  wire[45:0] T1986;
  wire[45:0] T1987;
  wire T1988;
  wire[46:0] twiddle3_1_49_imag;
  wire[46:0] T1989;
  wire[46:0] T1990;
  wire[46:0] T1991;
  wire[45:0] T1992;
  wire[45:0] T1993;
  wire T1994;
  wire T1995;
  wire[46:0] T1996;
  wire[46:0] twiddle3_1_50_imag;
  wire[46:0] T1997;
  wire[46:0] T1998;
  wire[46:0] T1999;
  wire[45:0] T2000;
  wire[45:0] T2001;
  wire T2002;
  wire[46:0] twiddle3_1_51_imag;
  wire[46:0] T2003;
  wire[46:0] T2004;
  wire[46:0] T2005;
  wire[44:0] T2006;
  wire[44:0] T2007;
  wire[1:0] T2008;
  wire T2009;
  wire T2010;
  wire T2011;
  wire[46:0] T2012;
  wire[46:0] T2013;
  wire[46:0] twiddle3_1_52_imag;
  wire[46:0] T2014;
  wire[46:0] T2015;
  wire[46:0] T2016;
  wire[44:0] T2017;
  wire[44:0] T2018;
  wire[1:0] T2019;
  wire T2020;
  wire[46:0] twiddle3_1_53_imag;
  wire[46:0] T2021;
  wire[46:0] T2022;
  wire[46:0] T2023;
  wire[44:0] T2024;
  wire[44:0] T2025;
  wire[1:0] T2026;
  wire T2027;
  wire T2028;
  wire[46:0] T2029;
  wire[46:0] twiddle3_1_54_imag;
  wire[46:0] T2030;
  wire[46:0] T2031;
  wire[46:0] T2032;
  wire[44:0] T2033;
  wire[44:0] T2034;
  wire[1:0] T2035;
  wire T2036;
  wire[46:0] twiddle3_1_55_imag;
  wire[46:0] T2037;
  wire[46:0] T2038;
  wire[46:0] T2039;
  wire[44:0] T2040;
  wire[44:0] T2041;
  wire[1:0] T2042;
  wire T2043;
  wire T2044;
  wire T2045;
  wire T2046;
  wire[46:0] T2047;
  wire[46:0] T2048;
  wire[46:0] T2049;
  wire[46:0] twiddle3_1_56_imag;
  wire[46:0] T2050;
  wire[46:0] T2051;
  wire[46:0] T2052;
  wire[43:0] T2053;
  wire[43:0] T2054;
  wire[2:0] T2055;
  wire T2056;
  wire[46:0] twiddle3_1_57_imag;
  wire[46:0] T2057;
  wire[46:0] T2058;
  wire[46:0] T2059;
  wire[43:0] T2060;
  wire[43:0] T2061;
  wire[2:0] T2062;
  wire T2063;
  wire T2064;
  wire[46:0] T2065;
  wire[46:0] twiddle3_1_58_imag;
  wire[46:0] T2066;
  wire[46:0] T2067;
  wire[46:0] T2068;
  wire[43:0] T2069;
  wire[43:0] T2070;
  wire[2:0] T2071;
  wire T2072;
  wire[46:0] twiddle3_1_59_imag;
  wire[46:0] T2073;
  wire[46:0] T2074;
  wire[46:0] T2075;
  wire[42:0] T2076;
  wire[42:0] T2077;
  wire[3:0] T2078;
  wire T2079;
  wire T2080;
  wire T2081;
  wire[46:0] T2082;
  wire[46:0] T2083;
  wire[46:0] twiddle3_1_60_imag;
  wire[46:0] T2084;
  wire[46:0] T2085;
  wire[46:0] T2086;
  wire[41:0] T2087;
  wire[41:0] T2088;
  wire[4:0] T2089;
  wire T2090;
  wire[46:0] twiddle3_1_61_imag;
  wire[46:0] T2091;
  wire[46:0] T2092;
  wire[46:0] T2093;
  wire[39:0] T2094;
  wire[39:0] T2095;
  wire[6:0] T2096;
  wire T2097;
  wire T2098;
  wire[46:0] T2099;
  wire[46:0] twiddle3_1_62_imag;
  wire[46:0] T2100;
  wire[46:0] T2101;
  wire[46:0] T2102;
  wire[42:0] T2103;
  wire[42:0] T2104;
  wire[3:0] T2105;
  wire T2106;
  wire[46:0] twiddle3_1_63_imag;
  wire[46:0] T2107;
  wire[46:0] T2108;
  wire[46:0] T2109;
  wire[42:0] T2110;
  wire[42:0] T2111;
  wire[3:0] T2112;
  wire T2113;
  wire T2114;
  wire T2115;
  wire T2116;
  wire T2117;
  wire T2118;
  wire T2119;
  wire T2120;
  wire[47:0] T2121;
  wire[46:0] T2122;
  wire[46:0] T2123;
  wire[46:0] T2124;
  wire[46:0] T2125;
  wire[46:0] T2126;
  wire[46:0] twiddle3_1_64_imag;
  wire[46:0] T2127;
  wire[46:0] T2128;
  wire[46:0] T2129;
  wire[43:0] T2130;
  wire[43:0] T2131;
  wire[2:0] T2132;
  wire T2133;
  wire[46:0] twiddle3_1_65_imag;
  wire[46:0] T2134;
  wire[46:0] T2135;
  wire[46:0] T2136;
  wire[43:0] T2137;
  wire[43:0] T2138;
  wire[2:0] T2139;
  wire T2140;
  wire T2141;
  wire[46:0] T2142;
  wire[46:0] twiddle3_1_66_imag;
  wire[46:0] T2143;
  wire[46:0] T2144;
  wire[46:0] T2145;
  wire[44:0] T2146;
  wire[44:0] T2147;
  wire[1:0] T2148;
  wire T2149;
  wire[46:0] twiddle3_1_67_imag;
  wire[46:0] T2150;
  wire[46:0] T2151;
  wire[46:0] T2152;
  wire[44:0] T2153;
  wire[44:0] T2154;
  wire[1:0] T2155;
  wire T2156;
  wire T2157;
  wire T2158;
  wire[46:0] T2159;
  wire[46:0] T2160;
  wire[46:0] twiddle3_1_68_imag;
  wire[46:0] T2161;
  wire[46:0] T2162;
  wire[46:0] T2163;
  wire[44:0] T2164;
  wire[44:0] T2165;
  wire[1:0] T2166;
  wire T2167;
  wire[46:0] twiddle3_1_69_imag;
  wire[46:0] T2168;
  wire[46:0] T2169;
  wire[46:0] T2170;
  wire[44:0] T2171;
  wire[44:0] T2172;
  wire[1:0] T2173;
  wire T2174;
  wire T2175;
  wire[46:0] T2176;
  wire[46:0] twiddle3_1_70_imag;
  wire[46:0] T2177;
  wire[46:0] T2178;
  wire[46:0] T2179;
  wire[44:0] T2180;
  wire[44:0] T2181;
  wire[1:0] T2182;
  wire T2183;
  wire[46:0] twiddle3_1_71_imag;
  wire[46:0] T2184;
  wire[46:0] T2185;
  wire[46:0] T2186;
  wire[45:0] T2187;
  wire[45:0] T2188;
  wire T2189;
  wire T2190;
  wire T2191;
  wire T2192;
  wire[46:0] T2193;
  wire[46:0] T2194;
  wire[46:0] T2195;
  wire[46:0] twiddle3_1_72_imag;
  wire[46:0] T2196;
  wire[46:0] T2197;
  wire[46:0] T2198;
  wire[45:0] T2199;
  wire[45:0] T2200;
  wire T2201;
  wire[46:0] twiddle3_1_73_imag;
  wire[46:0] T2202;
  wire[46:0] T2203;
  wire[46:0] T2204;
  wire[45:0] T2205;
  wire[45:0] T2206;
  wire T2207;
  wire T2208;
  wire[46:0] T2209;
  wire[46:0] twiddle3_1_74_imag;
  wire[46:0] T2210;
  wire[46:0] T2211;
  wire[46:0] T2212;
  wire[45:0] T2213;
  wire[45:0] T2214;
  wire T2215;
  wire[46:0] twiddle3_1_75_imag;
  wire[46:0] T2216;
  wire[46:0] T2217;
  wire[46:0] T2218;
  wire[45:0] T2219;
  wire[45:0] T2220;
  wire T2221;
  wire T2222;
  wire T2223;
  wire[46:0] T2224;
  wire[46:0] T2225;
  wire[46:0] twiddle3_1_76_imag;
  wire[46:0] T2226;
  wire[46:0] T2227;
  wire[46:0] T2228;
  wire[45:0] T2229;
  wire[45:0] T2230;
  wire T2231;
  wire[46:0] twiddle3_1_77_imag;
  wire[46:0] T2232;
  wire[46:0] T2233;
  wire[46:0] T2234;
  wire[45:0] T2235;
  wire[45:0] T2236;
  wire T2237;
  wire T2238;
  wire[46:0] T2239;
  wire[46:0] twiddle3_1_78_imag;
  wire[46:0] T2240;
  wire[46:0] T2241;
  wire[46:0] T2242;
  wire[45:0] T2243;
  wire[45:0] T2244;
  wire T2245;
  wire[46:0] twiddle3_1_79_imag;
  wire[46:0] T2246;
  wire[46:0] T2247;
  wire[46:0] T2248;
  wire[45:0] T2249;
  wire[45:0] T2250;
  wire T2251;
  wire T2252;
  wire T2253;
  wire T2254;
  wire T2255;
  wire[46:0] twiddle3_1_80_imag;
  wire[46:0] T2256;
  wire[46:0] T2257;
  wire[46:0] T2258;
  wire[45:0] T2259;
  wire[45:0] T2260;
  wire T2261;
  wire T2262;
  wire T2263;
  wire T2264;
  wire[15:0] T2265;
  wire[47:0] T2266;
  wire[47:0] T2267;
  wire[47:0] T2268;
  wire[47:0] T2269;
  wire[47:0] T2270;
  wire[47:0] T2271;
  wire[47:0] T2272;
  wire[47:0] twiddle3_1_0_real;
  wire[47:0] T2273;
  wire[16:0] T2274;
  wire[16:0] T2275;
  wire[30:0] T2276;
  wire T2277;
  wire[47:0] T2278;
  wire[47:0] T2279;
  wire[47:0] T2280;
  wire[46:0] twiddle3_1_1_real;
  wire[46:0] T2281;
  wire[41:0] T2282;
  wire[41:0] T2283;
  wire[4:0] T2284;
  wire T2285;
  wire[46:0] T2286;
  wire[46:0] T2287;
  wire T2288;
  wire T2289;
  wire[47:0] T2290;
  wire[46:0] T2291;
  wire[46:0] twiddle3_1_2_real;
  wire[46:0] T2292;
  wire[42:0] T2293;
  wire[42:0] T2294;
  wire[3:0] T2295;
  wire T2296;
  wire[46:0] T2297;
  wire[46:0] T2298;
  wire[46:0] twiddle3_1_3_real;
  wire[46:0] T2299;
  wire[43:0] T2300;
  wire[43:0] T2301;
  wire[2:0] T2302;
  wire T2303;
  wire[46:0] T2304;
  wire[46:0] T2305;
  wire T2306;
  wire T2307;
  wire T2308;
  wire[47:0] T2309;
  wire[46:0] T2310;
  wire[46:0] T2311;
  wire[46:0] twiddle3_1_4_real;
  wire[46:0] T2312;
  wire[43:0] T2313;
  wire[43:0] T2314;
  wire[2:0] T2315;
  wire T2316;
  wire[46:0] T2317;
  wire[46:0] T2318;
  wire[46:0] twiddle3_1_5_real;
  wire[46:0] T2319;
  wire[44:0] T2320;
  wire[44:0] T2321;
  wire[1:0] T2322;
  wire T2323;
  wire[46:0] T2324;
  wire[46:0] T2325;
  wire T2326;
  wire[46:0] T2327;
  wire[46:0] twiddle3_1_6_real;
  wire[46:0] T2328;
  wire[44:0] T2329;
  wire[44:0] T2330;
  wire[1:0] T2331;
  wire T2332;
  wire[46:0] T2333;
  wire[46:0] T2334;
  wire[46:0] twiddle3_1_7_real;
  wire[46:0] T2335;
  wire[44:0] T2336;
  wire[44:0] T2337;
  wire[1:0] T2338;
  wire T2339;
  wire[46:0] T2340;
  wire[46:0] T2341;
  wire T2342;
  wire T2343;
  wire T2344;
  wire T2345;
  wire[47:0] T2346;
  wire[46:0] T2347;
  wire[46:0] T2348;
  wire[46:0] T2349;
  wire[46:0] twiddle3_1_8_real;
  wire[46:0] T2350;
  wire[44:0] T2351;
  wire[44:0] T2352;
  wire[1:0] T2353;
  wire T2354;
  wire[46:0] T2355;
  wire[46:0] T2356;
  wire[46:0] twiddle3_1_9_real;
  wire[46:0] T2357;
  wire[44:0] T2358;
  wire[44:0] T2359;
  wire[1:0] T2360;
  wire T2361;
  wire[46:0] T2362;
  wire[46:0] T2363;
  wire T2364;
  wire[46:0] T2365;
  wire[46:0] twiddle3_1_10_real;
  wire[46:0] T2366;
  wire[45:0] T2367;
  wire[45:0] T2368;
  wire T2369;
  wire[46:0] T2370;
  wire[46:0] T2371;
  wire[46:0] twiddle3_1_11_real;
  wire[46:0] T2372;
  wire[45:0] T2373;
  wire[45:0] T2374;
  wire T2375;
  wire[46:0] T2376;
  wire[46:0] T2377;
  wire T2378;
  wire T2379;
  wire[46:0] T2380;
  wire[46:0] T2381;
  wire[46:0] twiddle3_1_12_real;
  wire[46:0] T2382;
  wire[45:0] T2383;
  wire[45:0] T2384;
  wire T2385;
  wire[46:0] T2386;
  wire[46:0] T2387;
  wire[46:0] twiddle3_1_13_real;
  wire[46:0] T2388;
  wire[45:0] T2389;
  wire[45:0] T2390;
  wire T2391;
  wire[46:0] T2392;
  wire[46:0] T2393;
  wire T2394;
  wire[46:0] T2395;
  wire[46:0] twiddle3_1_14_real;
  wire[46:0] T2396;
  wire[45:0] T2397;
  wire[45:0] T2398;
  wire T2399;
  wire[46:0] T2400;
  wire[46:0] T2401;
  wire[46:0] twiddle3_1_15_real;
  wire[46:0] T2402;
  wire[45:0] T2403;
  wire[45:0] T2404;
  wire T2405;
  wire[46:0] T2406;
  wire[46:0] T2407;
  wire T2408;
  wire T2409;
  wire T2410;
  wire T2411;
  wire T2412;
  wire[47:0] T2413;
  wire[46:0] T2414;
  wire[46:0] T2415;
  wire[46:0] T2416;
  wire[46:0] T2417;
  wire[46:0] twiddle3_1_16_real;
  wire[46:0] T2418;
  wire[45:0] T2419;
  wire[45:0] T2420;
  wire T2421;
  wire[46:0] T2422;
  wire[46:0] T2423;
  wire[46:0] twiddle3_1_17_real;
  wire[46:0] T2424;
  wire[45:0] T2425;
  wire[45:0] T2426;
  wire T2427;
  wire[46:0] T2428;
  wire[46:0] T2429;
  wire T2430;
  wire[46:0] T2431;
  wire[46:0] twiddle3_1_18_real;
  wire[46:0] T2432;
  wire[45:0] T2433;
  wire[45:0] T2434;
  wire T2435;
  wire[46:0] T2436;
  wire[46:0] T2437;
  wire[46:0] twiddle3_1_19_real;
  wire[46:0] T2438;
  wire[45:0] T2439;
  wire[45:0] T2440;
  wire T2441;
  wire[46:0] T2442;
  wire[46:0] T2443;
  wire T2444;
  wire T2445;
  wire[46:0] T2446;
  wire[46:0] T2447;
  wire[46:0] twiddle3_1_20_real;
  wire[46:0] T2448;
  wire[45:0] T2449;
  wire[45:0] T2450;
  wire T2451;
  wire[46:0] T2452;
  wire[46:0] T2453;
  wire[46:0] twiddle3_1_21_real;
  wire[46:0] T2454;
  wire[46:0] T2455;
  wire[46:0] T2456;
  wire[46:0] T2457;
  wire T2458;
  wire[46:0] T2459;
  wire[46:0] twiddle3_1_22_real;
  wire[46:0] T2460;
  wire[46:0] T2461;
  wire[46:0] T2462;
  wire[46:0] T2463;
  wire[46:0] twiddle3_1_23_real;
  wire[46:0] T2464;
  wire[46:0] T2465;
  wire[46:0] T2466;
  wire[46:0] T2467;
  wire T2468;
  wire T2469;
  wire T2470;
  wire[46:0] T2471;
  wire[46:0] T2472;
  wire[46:0] T2473;
  wire[46:0] twiddle3_1_24_real;
  wire[46:0] T2474;
  wire[46:0] T2475;
  wire[46:0] T2476;
  wire[46:0] T2477;
  wire[46:0] twiddle3_1_25_real;
  wire[46:0] T2478;
  wire[46:0] T2479;
  wire[46:0] T2480;
  wire[46:0] T2481;
  wire T2482;
  wire[46:0] T2483;
  wire[46:0] twiddle3_1_26_real;
  wire[46:0] T2484;
  wire[46:0] T2485;
  wire[46:0] T2486;
  wire[46:0] T2487;
  wire[46:0] twiddle3_1_27_real;
  wire[46:0] T2488;
  wire[46:0] T2489;
  wire[46:0] T2490;
  wire[46:0] T2491;
  wire T2492;
  wire T2493;
  wire[46:0] T2494;
  wire[46:0] T2495;
  wire[46:0] twiddle3_1_28_real;
  wire[46:0] T2496;
  wire[46:0] T2497;
  wire[46:0] T2498;
  wire[46:0] T2499;
  wire[46:0] twiddle3_1_29_real;
  wire[46:0] T2500;
  wire[46:0] T2501;
  wire[46:0] T2502;
  wire[46:0] T2503;
  wire T2504;
  wire[46:0] T2505;
  wire[46:0] twiddle3_1_30_real;
  wire[46:0] T2506;
  wire[46:0] T2507;
  wire[46:0] T2508;
  wire[46:0] T2509;
  wire[46:0] twiddle3_1_31_real;
  wire[46:0] T2510;
  wire[46:0] T2511;
  wire[46:0] T2512;
  wire[46:0] T2513;
  wire T2514;
  wire T2515;
  wire T2516;
  wire T2517;
  wire T2518;
  wire T2519;
  wire[47:0] T2520;
  wire[46:0] T2521;
  wire[46:0] T2522;
  wire[46:0] T2523;
  wire[46:0] T2524;
  wire[46:0] T2525;
  wire[46:0] twiddle3_1_32_real;
  wire[46:0] T2526;
  wire[46:0] T2527;
  wire[46:0] T2528;
  wire[46:0] T2529;
  wire[46:0] twiddle3_1_33_real;
  wire[46:0] T2530;
  wire[46:0] T2531;
  wire[46:0] T2532;
  wire[46:0] T2533;
  wire T2534;
  wire[46:0] T2535;
  wire[46:0] twiddle3_1_34_real;
  wire[46:0] T2536;
  wire[46:0] T2537;
  wire[46:0] T2538;
  wire[46:0] T2539;
  wire[46:0] twiddle3_1_35_real;
  wire[46:0] T2540;
  wire[46:0] T2541;
  wire[46:0] T2542;
  wire[46:0] T2543;
  wire T2544;
  wire T2545;
  wire[46:0] T2546;
  wire[46:0] T2547;
  wire[46:0] twiddle3_1_36_real;
  wire[46:0] T2548;
  wire[46:0] T2549;
  wire[46:0] T2550;
  wire[46:0] T2551;
  wire[46:0] twiddle3_1_37_real;
  wire[46:0] T2552;
  wire[46:0] T2553;
  wire[46:0] T2554;
  wire[46:0] T2555;
  wire T2556;
  wire[46:0] T2557;
  wire[46:0] twiddle3_1_38_real;
  wire[46:0] T2558;
  wire[46:0] T2559;
  wire[46:0] T2560;
  wire[46:0] T2561;
  wire[46:0] twiddle3_1_39_real;
  wire[46:0] T2562;
  wire[46:0] T2563;
  wire[46:0] T2564;
  wire[46:0] T2565;
  wire T2566;
  wire T2567;
  wire T2568;
  wire[46:0] T2569;
  wire[46:0] T2570;
  wire[46:0] T2571;
  wire[46:0] twiddle3_1_40_real;
  wire[46:0] T2572;
  wire[46:0] T2573;
  wire[46:0] T2574;
  wire[46:0] T2575;
  wire[46:0] twiddle3_1_41_real;
  wire[46:0] T2576;
  wire[46:0] T2577;
  wire[46:0] T2578;
  wire[45:0] T2579;
  wire[45:0] T2580;
  wire T2581;
  wire T2582;
  wire[46:0] T2583;
  wire[46:0] twiddle3_1_42_real;
  wire[46:0] T2584;
  wire[46:0] T2585;
  wire[46:0] T2586;
  wire[45:0] T2587;
  wire[45:0] T2588;
  wire T2589;
  wire[46:0] twiddle3_1_43_real;
  wire[46:0] T2590;
  wire[46:0] T2591;
  wire[46:0] T2592;
  wire[45:0] T2593;
  wire[45:0] T2594;
  wire T2595;
  wire T2596;
  wire T2597;
  wire[46:0] T2598;
  wire[46:0] T2599;
  wire[46:0] twiddle3_1_44_real;
  wire[46:0] T2600;
  wire[46:0] T2601;
  wire[46:0] T2602;
  wire[45:0] T2603;
  wire[45:0] T2604;
  wire T2605;
  wire[46:0] twiddle3_1_45_real;
  wire[46:0] T2606;
  wire[46:0] T2607;
  wire[46:0] T2608;
  wire[45:0] T2609;
  wire[45:0] T2610;
  wire T2611;
  wire T2612;
  wire[46:0] T2613;
  wire[46:0] twiddle3_1_46_real;
  wire[46:0] T2614;
  wire[46:0] T2615;
  wire[46:0] T2616;
  wire[45:0] T2617;
  wire[45:0] T2618;
  wire T2619;
  wire[46:0] twiddle3_1_47_real;
  wire[46:0] T2620;
  wire[46:0] T2621;
  wire[46:0] T2622;
  wire[45:0] T2623;
  wire[45:0] T2624;
  wire T2625;
  wire T2626;
  wire T2627;
  wire T2628;
  wire T2629;
  wire[46:0] T2630;
  wire[46:0] T2631;
  wire[46:0] T2632;
  wire[46:0] T2633;
  wire[46:0] twiddle3_1_48_real;
  wire[46:0] T2634;
  wire[46:0] T2635;
  wire[46:0] T2636;
  wire[45:0] T2637;
  wire[45:0] T2638;
  wire T2639;
  wire[46:0] twiddle3_1_49_real;
  wire[46:0] T2640;
  wire[46:0] T2641;
  wire[46:0] T2642;
  wire[45:0] T2643;
  wire[45:0] T2644;
  wire T2645;
  wire T2646;
  wire[46:0] T2647;
  wire[46:0] twiddle3_1_50_real;
  wire[46:0] T2648;
  wire[46:0] T2649;
  wire[46:0] T2650;
  wire[45:0] T2651;
  wire[45:0] T2652;
  wire T2653;
  wire[46:0] twiddle3_1_51_real;
  wire[46:0] T2654;
  wire[46:0] T2655;
  wire[46:0] T2656;
  wire[44:0] T2657;
  wire[44:0] T2658;
  wire[1:0] T2659;
  wire T2660;
  wire T2661;
  wire T2662;
  wire[46:0] T2663;
  wire[46:0] T2664;
  wire[46:0] twiddle3_1_52_real;
  wire[46:0] T2665;
  wire[46:0] T2666;
  wire[46:0] T2667;
  wire[44:0] T2668;
  wire[44:0] T2669;
  wire[1:0] T2670;
  wire T2671;
  wire[46:0] twiddle3_1_53_real;
  wire[46:0] T2672;
  wire[46:0] T2673;
  wire[46:0] T2674;
  wire[44:0] T2675;
  wire[44:0] T2676;
  wire[1:0] T2677;
  wire T2678;
  wire T2679;
  wire[46:0] T2680;
  wire[46:0] twiddle3_1_54_real;
  wire[46:0] T2681;
  wire[46:0] T2682;
  wire[46:0] T2683;
  wire[44:0] T2684;
  wire[44:0] T2685;
  wire[1:0] T2686;
  wire T2687;
  wire[46:0] twiddle3_1_55_real;
  wire[46:0] T2688;
  wire[46:0] T2689;
  wire[46:0] T2690;
  wire[44:0] T2691;
  wire[44:0] T2692;
  wire[1:0] T2693;
  wire T2694;
  wire T2695;
  wire T2696;
  wire T2697;
  wire[46:0] T2698;
  wire[46:0] T2699;
  wire[46:0] T2700;
  wire[46:0] twiddle3_1_56_real;
  wire[46:0] T2701;
  wire[46:0] T2702;
  wire[46:0] T2703;
  wire[43:0] T2704;
  wire[43:0] T2705;
  wire[2:0] T2706;
  wire T2707;
  wire[46:0] twiddle3_1_57_real;
  wire[46:0] T2708;
  wire[46:0] T2709;
  wire[46:0] T2710;
  wire[43:0] T2711;
  wire[43:0] T2712;
  wire[2:0] T2713;
  wire T2714;
  wire T2715;
  wire[46:0] T2716;
  wire[46:0] twiddle3_1_58_real;
  wire[46:0] T2717;
  wire[46:0] T2718;
  wire[46:0] T2719;
  wire[43:0] T2720;
  wire[43:0] T2721;
  wire[2:0] T2722;
  wire T2723;
  wire[46:0] twiddle3_1_59_real;
  wire[46:0] T2724;
  wire[46:0] T2725;
  wire[46:0] T2726;
  wire[42:0] T2727;
  wire[42:0] T2728;
  wire[3:0] T2729;
  wire T2730;
  wire T2731;
  wire T2732;
  wire[46:0] T2733;
  wire[46:0] T2734;
  wire[46:0] twiddle3_1_60_real;
  wire[46:0] T2735;
  wire[46:0] T2736;
  wire[46:0] T2737;
  wire[41:0] T2738;
  wire[41:0] T2739;
  wire[4:0] T2740;
  wire T2741;
  wire[46:0] twiddle3_1_61_real;
  wire[46:0] T2742;
  wire[46:0] T2743;
  wire[46:0] T2744;
  wire[39:0] T2745;
  wire[39:0] T2746;
  wire[6:0] T2747;
  wire T2748;
  wire T2749;
  wire[46:0] T2750;
  wire[46:0] twiddle3_1_62_real;
  wire[46:0] T2751;
  wire[46:0] T2752;
  wire[46:0] T2753;
  wire[42:0] T2754;
  wire[42:0] T2755;
  wire[3:0] T2756;
  wire T2757;
  wire[46:0] twiddle3_1_63_real;
  wire[46:0] T2758;
  wire[46:0] T2759;
  wire[46:0] T2760;
  wire[42:0] T2761;
  wire[42:0] T2762;
  wire[3:0] T2763;
  wire T2764;
  wire T2765;
  wire T2766;
  wire T2767;
  wire T2768;
  wire T2769;
  wire T2770;
  wire T2771;
  wire[47:0] T2772;
  wire[46:0] T2773;
  wire[46:0] T2774;
  wire[46:0] T2775;
  wire[46:0] T2776;
  wire[46:0] T2777;
  wire[46:0] twiddle3_1_64_real;
  wire[46:0] T2778;
  wire[46:0] T2779;
  wire[46:0] T2780;
  wire[43:0] T2781;
  wire[43:0] T2782;
  wire[2:0] T2783;
  wire T2784;
  wire[46:0] twiddle3_1_65_real;
  wire[46:0] T2785;
  wire[46:0] T2786;
  wire[46:0] T2787;
  wire[43:0] T2788;
  wire[43:0] T2789;
  wire[2:0] T2790;
  wire T2791;
  wire T2792;
  wire[46:0] T2793;
  wire[46:0] twiddle3_1_66_real;
  wire[46:0] T2794;
  wire[46:0] T2795;
  wire[46:0] T2796;
  wire[44:0] T2797;
  wire[44:0] T2798;
  wire[1:0] T2799;
  wire T2800;
  wire[46:0] twiddle3_1_67_real;
  wire[46:0] T2801;
  wire[46:0] T2802;
  wire[46:0] T2803;
  wire[44:0] T2804;
  wire[44:0] T2805;
  wire[1:0] T2806;
  wire T2807;
  wire T2808;
  wire T2809;
  wire[46:0] T2810;
  wire[46:0] T2811;
  wire[46:0] twiddle3_1_68_real;
  wire[46:0] T2812;
  wire[46:0] T2813;
  wire[46:0] T2814;
  wire[44:0] T2815;
  wire[44:0] T2816;
  wire[1:0] T2817;
  wire T2818;
  wire[46:0] twiddle3_1_69_real;
  wire[46:0] T2819;
  wire[46:0] T2820;
  wire[46:0] T2821;
  wire[44:0] T2822;
  wire[44:0] T2823;
  wire[1:0] T2824;
  wire T2825;
  wire T2826;
  wire[46:0] T2827;
  wire[46:0] twiddle3_1_70_real;
  wire[46:0] T2828;
  wire[46:0] T2829;
  wire[46:0] T2830;
  wire[44:0] T2831;
  wire[44:0] T2832;
  wire[1:0] T2833;
  wire T2834;
  wire[46:0] twiddle3_1_71_real;
  wire[46:0] T2835;
  wire[46:0] T2836;
  wire[46:0] T2837;
  wire[45:0] T2838;
  wire[45:0] T2839;
  wire T2840;
  wire T2841;
  wire T2842;
  wire T2843;
  wire[46:0] T2844;
  wire[46:0] T2845;
  wire[46:0] T2846;
  wire[46:0] twiddle3_1_72_real;
  wire[46:0] T2847;
  wire[46:0] T2848;
  wire[46:0] T2849;
  wire[45:0] T2850;
  wire[45:0] T2851;
  wire T2852;
  wire[46:0] twiddle3_1_73_real;
  wire[46:0] T2853;
  wire[46:0] T2854;
  wire[46:0] T2855;
  wire[45:0] T2856;
  wire[45:0] T2857;
  wire T2858;
  wire T2859;
  wire[46:0] T2860;
  wire[46:0] twiddle3_1_74_real;
  wire[46:0] T2861;
  wire[46:0] T2862;
  wire[46:0] T2863;
  wire[45:0] T2864;
  wire[45:0] T2865;
  wire T2866;
  wire[46:0] twiddle3_1_75_real;
  wire[46:0] T2867;
  wire[46:0] T2868;
  wire[46:0] T2869;
  wire[45:0] T2870;
  wire[45:0] T2871;
  wire T2872;
  wire T2873;
  wire T2874;
  wire[46:0] T2875;
  wire[46:0] T2876;
  wire[46:0] twiddle3_1_76_real;
  wire[46:0] T2877;
  wire[46:0] T2878;
  wire[46:0] T2879;
  wire[45:0] T2880;
  wire[45:0] T2881;
  wire T2882;
  wire[46:0] twiddle3_1_77_real;
  wire[46:0] T2883;
  wire[46:0] T2884;
  wire[46:0] T2885;
  wire[45:0] T2886;
  wire[45:0] T2887;
  wire T2888;
  wire T2889;
  wire[46:0] T2890;
  wire[46:0] twiddle3_1_78_real;
  wire[46:0] T2891;
  wire[46:0] T2892;
  wire[46:0] T2893;
  wire[45:0] T2894;
  wire[45:0] T2895;
  wire T2896;
  wire[46:0] twiddle3_1_79_real;
  wire[46:0] T2897;
  wire[46:0] T2898;
  wire[46:0] T2899;
  wire[45:0] T2900;
  wire[45:0] T2901;
  wire T2902;
  wire T2903;
  wire T2904;
  wire T2905;
  wire T2906;
  wire[46:0] twiddle3_1_80_real;
  wire[46:0] T2907;
  wire[46:0] T2908;
  wire[46:0] T2909;
  wire[45:0] T2910;
  wire[45:0] T2911;
  wire T2912;
  wire T2913;
  wire T2914;
  wire T2915;
  wire[15:0] T2916;
  wire[47:0] T2917;
  wire[47:0] T2918;
  wire[47:0] T2919;
  wire[47:0] T2920;
  wire[47:0] T2921;
  wire[47:0] T2922;
  wire[47:0] T2923;
  wire[47:0] T2924;
  wire[47:0] T2925;
  wire[47:0] twiddle4_3_0_imag;
  wire[47:0] T2926;
  wire[16:0] T2927;
  wire[16:0] T2928;
  wire[30:0] T2929;
  wire T2930;
  wire[47:0] T2931;
  wire[47:0] T2932;
  wire[47:0] T2933;
  wire[46:0] twiddle4_3_1_imag;
  wire[46:0] T2934;
  wire[40:0] T2935;
  wire[40:0] T2936;
  wire[5:0] T2937;
  wire T2938;
  wire[46:0] T2939;
  wire[46:0] T2940;
  wire T2941;
  wire T2942;
  wire[8:0] T2943;
  wire[8:0] T2944;
  wire[47:0] T2945;
  wire[46:0] T2946;
  wire[46:0] twiddle4_3_2_imag;
  wire[46:0] T2947;
  wire[41:0] T2948;
  wire[41:0] T2949;
  wire[4:0] T2950;
  wire T2951;
  wire[46:0] T2952;
  wire[46:0] T2953;
  wire[46:0] twiddle4_3_3_imag;
  wire[46:0] T2954;
  wire[41:0] T2955;
  wire[41:0] T2956;
  wire[4:0] T2957;
  wire T2958;
  wire[46:0] T2959;
  wire[46:0] T2960;
  wire T2961;
  wire T2962;
  wire T2963;
  wire[47:0] T2964;
  wire[46:0] T2965;
  wire[46:0] T2966;
  wire[46:0] twiddle4_3_4_imag;
  wire[46:0] T2967;
  wire[42:0] T2968;
  wire[42:0] T2969;
  wire[3:0] T2970;
  wire T2971;
  wire[46:0] T2972;
  wire[46:0] T2973;
  wire[46:0] twiddle4_3_5_imag;
  wire[46:0] T2974;
  wire[42:0] T2975;
  wire[42:0] T2976;
  wire[3:0] T2977;
  wire T2978;
  wire[46:0] T2979;
  wire[46:0] T2980;
  wire T2981;
  wire[46:0] T2982;
  wire[46:0] twiddle4_3_6_imag;
  wire[46:0] T2983;
  wire[42:0] T2984;
  wire[42:0] T2985;
  wire[3:0] T2986;
  wire T2987;
  wire[46:0] T2988;
  wire[46:0] T2989;
  wire[46:0] twiddle4_3_7_imag;
  wire[46:0] T2990;
  wire[43:0] T2991;
  wire[43:0] T2992;
  wire[2:0] T2993;
  wire T2994;
  wire[46:0] T2995;
  wire[46:0] T2996;
  wire T2997;
  wire T2998;
  wire T2999;
  wire T3000;
  wire[47:0] T3001;
  wire[46:0] T3002;
  wire[46:0] T3003;
  wire[46:0] T3004;
  wire[46:0] twiddle4_3_8_imag;
  wire[46:0] T3005;
  wire[43:0] T3006;
  wire[43:0] T3007;
  wire[2:0] T3008;
  wire T3009;
  wire[46:0] T3010;
  wire[46:0] T3011;
  wire[46:0] twiddle4_3_9_imag;
  wire[46:0] T3012;
  wire[43:0] T3013;
  wire[43:0] T3014;
  wire[2:0] T3015;
  wire T3016;
  wire[46:0] T3017;
  wire[46:0] T3018;
  wire T3019;
  wire[46:0] T3020;
  wire[46:0] twiddle4_3_10_imag;
  wire[46:0] T3021;
  wire[43:0] T3022;
  wire[43:0] T3023;
  wire[2:0] T3024;
  wire T3025;
  wire[46:0] T3026;
  wire[46:0] T3027;
  wire[46:0] twiddle4_3_11_imag;
  wire[46:0] T3028;
  wire[43:0] T3029;
  wire[43:0] T3030;
  wire[2:0] T3031;
  wire T3032;
  wire[46:0] T3033;
  wire[46:0] T3034;
  wire T3035;
  wire T3036;
  wire[46:0] T3037;
  wire[46:0] T3038;
  wire[46:0] twiddle4_3_12_imag;
  wire[46:0] T3039;
  wire[43:0] T3040;
  wire[43:0] T3041;
  wire[2:0] T3042;
  wire T3043;
  wire[46:0] T3044;
  wire[46:0] T3045;
  wire[46:0] twiddle4_3_13_imag;
  wire[46:0] T3046;
  wire[43:0] T3047;
  wire[43:0] T3048;
  wire[2:0] T3049;
  wire T3050;
  wire[46:0] T3051;
  wire[46:0] T3052;
  wire T3053;
  wire[46:0] T3054;
  wire[46:0] twiddle4_3_14_imag;
  wire[46:0] T3055;
  wire[44:0] T3056;
  wire[44:0] T3057;
  wire[1:0] T3058;
  wire T3059;
  wire[46:0] T3060;
  wire[46:0] T3061;
  wire[46:0] twiddle4_3_15_imag;
  wire[46:0] T3062;
  wire[44:0] T3063;
  wire[44:0] T3064;
  wire[1:0] T3065;
  wire T3066;
  wire[46:0] T3067;
  wire[46:0] T3068;
  wire T3069;
  wire T3070;
  wire T3071;
  wire T3072;
  wire T3073;
  wire[47:0] T3074;
  wire[46:0] T3075;
  wire[46:0] T3076;
  wire[46:0] T3077;
  wire[46:0] T3078;
  wire[46:0] twiddle4_3_16_imag;
  wire[46:0] T3079;
  wire[44:0] T3080;
  wire[44:0] T3081;
  wire[1:0] T3082;
  wire T3083;
  wire[46:0] T3084;
  wire[46:0] T3085;
  wire[46:0] twiddle4_3_17_imag;
  wire[46:0] T3086;
  wire[44:0] T3087;
  wire[44:0] T3088;
  wire[1:0] T3089;
  wire T3090;
  wire[46:0] T3091;
  wire[46:0] T3092;
  wire T3093;
  wire[46:0] T3094;
  wire[46:0] twiddle4_3_18_imag;
  wire[46:0] T3095;
  wire[44:0] T3096;
  wire[44:0] T3097;
  wire[1:0] T3098;
  wire T3099;
  wire[46:0] T3100;
  wire[46:0] T3101;
  wire[46:0] twiddle4_3_19_imag;
  wire[46:0] T3102;
  wire[44:0] T3103;
  wire[44:0] T3104;
  wire[1:0] T3105;
  wire T3106;
  wire[46:0] T3107;
  wire[46:0] T3108;
  wire T3109;
  wire T3110;
  wire[46:0] T3111;
  wire[46:0] T3112;
  wire[46:0] twiddle4_3_20_imag;
  wire[46:0] T3113;
  wire[44:0] T3114;
  wire[44:0] T3115;
  wire[1:0] T3116;
  wire T3117;
  wire[46:0] T3118;
  wire[46:0] T3119;
  wire[46:0] twiddle4_3_21_imag;
  wire[46:0] T3120;
  wire[44:0] T3121;
  wire[44:0] T3122;
  wire[1:0] T3123;
  wire T3124;
  wire[46:0] T3125;
  wire[46:0] T3126;
  wire T3127;
  wire[46:0] T3128;
  wire[46:0] twiddle4_3_22_imag;
  wire[46:0] T3129;
  wire[44:0] T3130;
  wire[44:0] T3131;
  wire[1:0] T3132;
  wire T3133;
  wire[46:0] T3134;
  wire[46:0] T3135;
  wire[46:0] twiddle4_3_23_imag;
  wire[46:0] T3136;
  wire[44:0] T3137;
  wire[44:0] T3138;
  wire[1:0] T3139;
  wire T3140;
  wire[46:0] T3141;
  wire[46:0] T3142;
  wire T3143;
  wire T3144;
  wire T3145;
  wire[46:0] T3146;
  wire[46:0] T3147;
  wire[46:0] T3148;
  wire[46:0] twiddle4_3_24_imag;
  wire[46:0] T3149;
  wire[44:0] T3150;
  wire[44:0] T3151;
  wire[1:0] T3152;
  wire T3153;
  wire[46:0] T3154;
  wire[46:0] T3155;
  wire[46:0] twiddle4_3_25_imag;
  wire[46:0] T3156;
  wire[44:0] T3157;
  wire[44:0] T3158;
  wire[1:0] T3159;
  wire T3160;
  wire[46:0] T3161;
  wire[46:0] T3162;
  wire T3163;
  wire[46:0] T3164;
  wire[46:0] twiddle4_3_26_imag;
  wire[46:0] T3165;
  wire[44:0] T3166;
  wire[44:0] T3167;
  wire[1:0] T3168;
  wire T3169;
  wire[46:0] T3170;
  wire[46:0] T3171;
  wire[46:0] twiddle4_3_27_imag;
  wire[46:0] T3172;
  wire[44:0] T3173;
  wire[44:0] T3174;
  wire[1:0] T3175;
  wire T3176;
  wire[46:0] T3177;
  wire[46:0] T3178;
  wire T3179;
  wire T3180;
  wire[46:0] T3181;
  wire[46:0] T3182;
  wire[46:0] twiddle4_3_28_imag;
  wire[46:0] T3183;
  wire[45:0] T3184;
  wire[45:0] T3185;
  wire T3186;
  wire[46:0] T3187;
  wire[46:0] T3188;
  wire[46:0] twiddle4_3_29_imag;
  wire[46:0] T3189;
  wire[45:0] T3190;
  wire[45:0] T3191;
  wire T3192;
  wire[46:0] T3193;
  wire[46:0] T3194;
  wire T3195;
  wire[46:0] T3196;
  wire[46:0] twiddle4_3_30_imag;
  wire[46:0] T3197;
  wire[45:0] T3198;
  wire[45:0] T3199;
  wire T3200;
  wire[46:0] T3201;
  wire[46:0] T3202;
  wire[46:0] twiddle4_3_31_imag;
  wire[46:0] T3203;
  wire[45:0] T3204;
  wire[45:0] T3205;
  wire T3206;
  wire[46:0] T3207;
  wire[46:0] T3208;
  wire T3209;
  wire T3210;
  wire T3211;
  wire T3212;
  wire T3213;
  wire T3214;
  wire[47:0] T3215;
  wire[46:0] T3216;
  wire[46:0] T3217;
  wire[46:0] T3218;
  wire[46:0] T3219;
  wire[46:0] T3220;
  wire[46:0] twiddle4_3_32_imag;
  wire[46:0] T3221;
  wire[45:0] T3222;
  wire[45:0] T3223;
  wire T3224;
  wire[46:0] T3225;
  wire[46:0] T3226;
  wire[46:0] twiddle4_3_33_imag;
  wire[46:0] T3227;
  wire[45:0] T3228;
  wire[45:0] T3229;
  wire T3230;
  wire[46:0] T3231;
  wire[46:0] T3232;
  wire T3233;
  wire[46:0] T3234;
  wire[46:0] twiddle4_3_34_imag;
  wire[46:0] T3235;
  wire[45:0] T3236;
  wire[45:0] T3237;
  wire T3238;
  wire[46:0] T3239;
  wire[46:0] T3240;
  wire[46:0] twiddle4_3_35_imag;
  wire[46:0] T3241;
  wire[45:0] T3242;
  wire[45:0] T3243;
  wire T3244;
  wire[46:0] T3245;
  wire[46:0] T3246;
  wire T3247;
  wire T3248;
  wire[46:0] T3249;
  wire[46:0] T3250;
  wire[46:0] twiddle4_3_36_imag;
  wire[46:0] T3251;
  wire[45:0] T3252;
  wire[45:0] T3253;
  wire T3254;
  wire[46:0] T3255;
  wire[46:0] T3256;
  wire[46:0] twiddle4_3_37_imag;
  wire[46:0] T3257;
  wire[45:0] T3258;
  wire[45:0] T3259;
  wire T3260;
  wire[46:0] T3261;
  wire[46:0] T3262;
  wire T3263;
  wire[46:0] T3264;
  wire[46:0] twiddle4_3_38_imag;
  wire[46:0] T3265;
  wire[45:0] T3266;
  wire[45:0] T3267;
  wire T3268;
  wire[46:0] T3269;
  wire[46:0] T3270;
  wire[46:0] twiddle4_3_39_imag;
  wire[46:0] T3271;
  wire[45:0] T3272;
  wire[45:0] T3273;
  wire T3274;
  wire[46:0] T3275;
  wire[46:0] T3276;
  wire T3277;
  wire T3278;
  wire T3279;
  wire[46:0] T3280;
  wire[46:0] T3281;
  wire[46:0] T3282;
  wire[46:0] twiddle4_3_40_imag;
  wire[46:0] T3283;
  wire[45:0] T3284;
  wire[45:0] T3285;
  wire T3286;
  wire[46:0] T3287;
  wire[46:0] T3288;
  wire[46:0] twiddle4_3_41_imag;
  wire[46:0] T3289;
  wire[45:0] T3290;
  wire[45:0] T3291;
  wire T3292;
  wire[46:0] T3293;
  wire[46:0] T3294;
  wire T3295;
  wire[46:0] T3296;
  wire[46:0] twiddle4_3_42_imag;
  wire[46:0] T3297;
  wire[45:0] T3298;
  wire[45:0] T3299;
  wire T3300;
  wire[46:0] T3301;
  wire[46:0] T3302;
  wire[46:0] twiddle4_3_43_imag;
  wire[46:0] T3303;
  wire[45:0] T3304;
  wire[45:0] T3305;
  wire T3306;
  wire[46:0] T3307;
  wire[46:0] T3308;
  wire T3309;
  wire T3310;
  wire[46:0] T3311;
  wire[46:0] T3312;
  wire[46:0] twiddle4_3_44_imag;
  wire[46:0] T3313;
  wire[45:0] T3314;
  wire[45:0] T3315;
  wire T3316;
  wire[46:0] T3317;
  wire[46:0] T3318;
  wire[46:0] twiddle4_3_45_imag;
  wire[46:0] T3319;
  wire[45:0] T3320;
  wire[45:0] T3321;
  wire T3322;
  wire[46:0] T3323;
  wire[46:0] T3324;
  wire T3325;
  wire[46:0] T3326;
  wire[46:0] twiddle4_3_46_imag;
  wire[46:0] T3327;
  wire[45:0] T3328;
  wire[45:0] T3329;
  wire T3330;
  wire[46:0] T3331;
  wire[46:0] T3332;
  wire[46:0] twiddle4_3_47_imag;
  wire[46:0] T3333;
  wire[45:0] T3334;
  wire[45:0] T3335;
  wire T3336;
  wire[46:0] T3337;
  wire[46:0] T3338;
  wire T3339;
  wire T3340;
  wire T3341;
  wire T3342;
  wire[46:0] T3343;
  wire[46:0] T3344;
  wire[46:0] T3345;
  wire[46:0] T3346;
  wire[46:0] twiddle4_3_48_imag;
  wire[46:0] T3347;
  wire[45:0] T3348;
  wire[45:0] T3349;
  wire T3350;
  wire[46:0] T3351;
  wire[46:0] T3352;
  wire[46:0] twiddle4_3_49_imag;
  wire[46:0] T3353;
  wire[45:0] T3354;
  wire[45:0] T3355;
  wire T3356;
  wire[46:0] T3357;
  wire[46:0] T3358;
  wire T3359;
  wire[46:0] T3360;
  wire[46:0] twiddle4_3_50_imag;
  wire[46:0] T3361;
  wire[45:0] T3362;
  wire[45:0] T3363;
  wire T3364;
  wire[46:0] T3365;
  wire[46:0] T3366;
  wire[46:0] twiddle4_3_51_imag;
  wire[46:0] T3367;
  wire[45:0] T3368;
  wire[45:0] T3369;
  wire T3370;
  wire[46:0] T3371;
  wire[46:0] T3372;
  wire T3373;
  wire T3374;
  wire[46:0] T3375;
  wire[46:0] T3376;
  wire[46:0] twiddle4_3_52_imag;
  wire[46:0] T3377;
  wire[45:0] T3378;
  wire[45:0] T3379;
  wire T3380;
  wire[46:0] T3381;
  wire[46:0] T3382;
  wire[46:0] twiddle4_3_53_imag;
  wire[46:0] T3383;
  wire[45:0] T3384;
  wire[45:0] T3385;
  wire T3386;
  wire[46:0] T3387;
  wire[46:0] T3388;
  wire T3389;
  wire[46:0] T3390;
  wire[46:0] twiddle4_3_54_imag;
  wire[46:0] T3391;
  wire[45:0] T3392;
  wire[45:0] T3393;
  wire T3394;
  wire[46:0] T3395;
  wire[46:0] T3396;
  wire[46:0] twiddle4_3_55_imag;
  wire[46:0] T3397;
  wire[45:0] T3398;
  wire[45:0] T3399;
  wire T3400;
  wire[46:0] T3401;
  wire[46:0] T3402;
  wire T3403;
  wire T3404;
  wire T3405;
  wire[46:0] T3406;
  wire[46:0] T3407;
  wire[46:0] T3408;
  wire[46:0] twiddle4_3_56_imag;
  wire[46:0] T3409;
  wire[45:0] T3410;
  wire[45:0] T3411;
  wire T3412;
  wire[46:0] T3413;
  wire[46:0] T3414;
  wire[46:0] twiddle4_3_57_imag;
  wire[46:0] T3415;
  wire[46:0] T3416;
  wire[46:0] T3417;
  wire[46:0] T3418;
  wire T3419;
  wire[46:0] T3420;
  wire[46:0] twiddle4_3_58_imag;
  wire[46:0] T3421;
  wire[46:0] T3422;
  wire[46:0] T3423;
  wire[46:0] T3424;
  wire[46:0] twiddle4_3_59_imag;
  wire[46:0] T3425;
  wire[46:0] T3426;
  wire[46:0] T3427;
  wire[46:0] T3428;
  wire T3429;
  wire T3430;
  wire[46:0] T3431;
  wire[46:0] T3432;
  wire[46:0] twiddle4_3_60_imag;
  wire[46:0] T3433;
  wire[46:0] T3434;
  wire[46:0] T3435;
  wire[46:0] T3436;
  wire[46:0] twiddle4_3_61_imag;
  wire[46:0] T3437;
  wire[46:0] T3438;
  wire[46:0] T3439;
  wire[46:0] T3440;
  wire T3441;
  wire[46:0] T3442;
  wire[46:0] twiddle4_3_62_imag;
  wire[46:0] T3443;
  wire[46:0] T3444;
  wire[46:0] T3445;
  wire[46:0] T3446;
  wire[46:0] twiddle4_3_63_imag;
  wire[46:0] T3447;
  wire[46:0] T3448;
  wire[46:0] T3449;
  wire[46:0] T3450;
  wire T3451;
  wire T3452;
  wire T3453;
  wire T3454;
  wire T3455;
  wire T3456;
  wire T3457;
  wire[47:0] T3458;
  wire[46:0] T3459;
  wire[46:0] T3460;
  wire[46:0] T3461;
  wire[46:0] T3462;
  wire[46:0] T3463;
  wire[46:0] T3464;
  wire[46:0] twiddle4_3_64_imag;
  wire[46:0] T3465;
  wire[46:0] T3466;
  wire[46:0] T3467;
  wire[46:0] T3468;
  wire[46:0] twiddle4_3_65_imag;
  wire[46:0] T3469;
  wire[46:0] T3470;
  wire[46:0] T3471;
  wire[46:0] T3472;
  wire T3473;
  wire[46:0] T3474;
  wire[46:0] twiddle4_3_66_imag;
  wire[46:0] T3475;
  wire[46:0] T3476;
  wire[46:0] T3477;
  wire[46:0] T3478;
  wire[46:0] twiddle4_3_67_imag;
  wire[46:0] T3479;
  wire[46:0] T3480;
  wire[46:0] T3481;
  wire[46:0] T3482;
  wire T3483;
  wire T3484;
  wire[46:0] T3485;
  wire[46:0] T3486;
  wire[46:0] twiddle4_3_68_imag;
  wire[46:0] T3487;
  wire[46:0] T3488;
  wire[46:0] T3489;
  wire[46:0] T3490;
  wire[46:0] twiddle4_3_69_imag;
  wire[46:0] T3491;
  wire[46:0] T3492;
  wire[46:0] T3493;
  wire[46:0] T3494;
  wire T3495;
  wire[46:0] T3496;
  wire[46:0] twiddle4_3_70_imag;
  wire[46:0] T3497;
  wire[46:0] T3498;
  wire[46:0] T3499;
  wire[46:0] T3500;
  wire[46:0] twiddle4_3_71_imag;
  wire[46:0] T3501;
  wire[46:0] T3502;
  wire[46:0] T3503;
  wire[46:0] T3504;
  wire T3505;
  wire T3506;
  wire T3507;
  wire[46:0] T3508;
  wire[46:0] T3509;
  wire[46:0] T3510;
  wire[46:0] twiddle4_3_72_imag;
  wire[46:0] T3511;
  wire[46:0] T3512;
  wire[46:0] T3513;
  wire[46:0] T3514;
  wire[46:0] twiddle4_3_73_imag;
  wire[46:0] T3515;
  wire[46:0] T3516;
  wire[46:0] T3517;
  wire[46:0] T3518;
  wire T3519;
  wire[46:0] T3520;
  wire[46:0] twiddle4_3_74_imag;
  wire[46:0] T3521;
  wire[46:0] T3522;
  wire[46:0] T3523;
  wire[46:0] T3524;
  wire[46:0] twiddle4_3_75_imag;
  wire[46:0] T3525;
  wire[46:0] T3526;
  wire[46:0] T3527;
  wire[46:0] T3528;
  wire T3529;
  wire T3530;
  wire[46:0] T3531;
  wire[46:0] T3532;
  wire[46:0] twiddle4_3_76_imag;
  wire[46:0] T3533;
  wire[46:0] T3534;
  wire[46:0] T3535;
  wire[46:0] T3536;
  wire[46:0] twiddle4_3_77_imag;
  wire[46:0] T3537;
  wire[46:0] T3538;
  wire[46:0] T3539;
  wire[46:0] T3540;
  wire T3541;
  wire[46:0] T3542;
  wire[46:0] twiddle4_3_78_imag;
  wire[46:0] T3543;
  wire[46:0] T3544;
  wire[46:0] T3545;
  wire[46:0] T3546;
  wire[46:0] twiddle4_3_79_imag;
  wire[46:0] T3547;
  wire[46:0] T3548;
  wire[46:0] T3549;
  wire[46:0] T3550;
  wire T3551;
  wire T3552;
  wire T3553;
  wire T3554;
  wire[46:0] T3555;
  wire[46:0] T3556;
  wire[46:0] T3557;
  wire[46:0] T3558;
  wire[46:0] twiddle4_3_80_imag;
  wire[46:0] T3559;
  wire[46:0] T3560;
  wire[46:0] T3561;
  wire[46:0] T3562;
  wire[46:0] twiddle4_3_81_imag;
  wire[46:0] T3563;
  wire[46:0] T3564;
  wire[46:0] T3565;
  wire[46:0] T3566;
  wire T3567;
  wire[46:0] T3568;
  wire[46:0] twiddle4_3_82_imag;
  wire[46:0] T3569;
  wire[46:0] T3570;
  wire[46:0] T3571;
  wire[46:0] T3572;
  wire[46:0] twiddle4_3_83_imag;
  wire[46:0] T3573;
  wire[46:0] T3574;
  wire[46:0] T3575;
  wire[46:0] T3576;
  wire T3577;
  wire T3578;
  wire[46:0] T3579;
  wire[46:0] T3580;
  wire[46:0] twiddle4_3_84_imag;
  wire[46:0] T3581;
  wire[46:0] T3582;
  wire[46:0] T3583;
  wire[46:0] T3584;
  wire[46:0] twiddle4_3_85_imag;
  wire[46:0] T3585;
  wire[46:0] T3586;
  wire[46:0] T3587;
  wire[46:0] T3588;
  wire T3589;
  wire[46:0] T3590;
  wire[46:0] twiddle4_3_86_imag;
  wire[46:0] T3591;
  wire[46:0] T3592;
  wire[46:0] T3593;
  wire[46:0] T3594;
  wire[46:0] twiddle4_3_87_imag;
  wire[46:0] T3595;
  wire[46:0] T3596;
  wire[46:0] T3597;
  wire[46:0] T3598;
  wire T3599;
  wire T3600;
  wire T3601;
  wire[46:0] T3602;
  wire[46:0] T3603;
  wire[46:0] T3604;
  wire[46:0] twiddle4_3_88_imag;
  wire[46:0] T3605;
  wire[46:0] T3606;
  wire[46:0] T3607;
  wire[46:0] T3608;
  wire[46:0] twiddle4_3_89_imag;
  wire[46:0] T3609;
  wire[46:0] T3610;
  wire[46:0] T3611;
  wire[46:0] T3612;
  wire T3613;
  wire[46:0] T3614;
  wire[46:0] twiddle4_3_90_imag;
  wire[46:0] T3615;
  wire[46:0] T3616;
  wire[46:0] T3617;
  wire[46:0] T3618;
  wire[46:0] twiddle4_3_91_imag;
  wire[46:0] T3619;
  wire[46:0] T3620;
  wire[46:0] T3621;
  wire[46:0] T3622;
  wire T3623;
  wire T3624;
  wire[46:0] T3625;
  wire[46:0] T3626;
  wire[46:0] twiddle4_3_92_imag;
  wire[46:0] T3627;
  wire[46:0] T3628;
  wire[46:0] T3629;
  wire[46:0] T3630;
  wire[46:0] twiddle4_3_93_imag;
  wire[46:0] T3631;
  wire[46:0] T3632;
  wire[46:0] T3633;
  wire[46:0] T3634;
  wire T3635;
  wire[46:0] T3636;
  wire[46:0] twiddle4_3_94_imag;
  wire[46:0] T3637;
  wire[46:0] T3638;
  wire[46:0] T3639;
  wire[46:0] T3640;
  wire[46:0] twiddle4_3_95_imag;
  wire[46:0] T3641;
  wire[46:0] T3642;
  wire[46:0] T3643;
  wire[46:0] T3644;
  wire T3645;
  wire T3646;
  wire T3647;
  wire T3648;
  wire T3649;
  wire[46:0] T3650;
  wire[46:0] T3651;
  wire[46:0] T3652;
  wire[46:0] T3653;
  wire[46:0] T3654;
  wire[46:0] twiddle4_3_96_imag;
  wire[46:0] T3655;
  wire[46:0] T3656;
  wire[46:0] T3657;
  wire[46:0] T3658;
  wire[46:0] twiddle4_3_97_imag;
  wire[46:0] T3659;
  wire[46:0] T3660;
  wire[46:0] T3661;
  wire[46:0] T3662;
  wire T3663;
  wire[46:0] T3664;
  wire[46:0] twiddle4_3_98_imag;
  wire[46:0] T3665;
  wire[46:0] T3666;
  wire[46:0] T3667;
  wire[46:0] T3668;
  wire[46:0] twiddle4_3_99_imag;
  wire[46:0] T3669;
  wire[46:0] T3670;
  wire[46:0] T3671;
  wire[46:0] T3672;
  wire T3673;
  wire T3674;
  wire[46:0] T3675;
  wire[46:0] T3676;
  wire[46:0] twiddle4_3_100_imag;
  wire[46:0] T3677;
  wire[46:0] T3678;
  wire[46:0] T3679;
  wire[46:0] T3680;
  wire[46:0] twiddle4_3_101_imag;
  wire[46:0] T3681;
  wire[46:0] T3682;
  wire[46:0] T3683;
  wire[46:0] T3684;
  wire T3685;
  wire[46:0] T3686;
  wire[46:0] twiddle4_3_102_imag;
  wire[46:0] T3687;
  wire[46:0] T3688;
  wire[46:0] T3689;
  wire[46:0] T3690;
  wire[46:0] twiddle4_3_103_imag;
  wire[46:0] T3691;
  wire[46:0] T3692;
  wire[46:0] T3693;
  wire[46:0] T3694;
  wire T3695;
  wire T3696;
  wire T3697;
  wire[46:0] T3698;
  wire[46:0] T3699;
  wire[46:0] T3700;
  wire[46:0] twiddle4_3_104_imag;
  wire[46:0] T3701;
  wire[46:0] T3702;
  wire[46:0] T3703;
  wire[46:0] T3704;
  wire[46:0] twiddle4_3_105_imag;
  wire[46:0] T3705;
  wire[46:0] T3706;
  wire[46:0] T3707;
  wire[46:0] T3708;
  wire T3709;
  wire[46:0] T3710;
  wire[46:0] twiddle4_3_106_imag;
  wire[46:0] T3711;
  wire[46:0] T3712;
  wire[46:0] T3713;
  wire[46:0] T3714;
  wire[46:0] twiddle4_3_107_imag;
  wire[46:0] T3715;
  wire[46:0] T3716;
  wire[46:0] T3717;
  wire[46:0] T3718;
  wire T3719;
  wire T3720;
  wire[46:0] T3721;
  wire[46:0] T3722;
  wire[46:0] twiddle4_3_108_imag;
  wire[46:0] T3723;
  wire[46:0] T3724;
  wire[46:0] T3725;
  wire[46:0] T3726;
  wire[46:0] twiddle4_3_109_imag;
  wire[46:0] T3727;
  wire[46:0] T3728;
  wire[46:0] T3729;
  wire[46:0] T3730;
  wire T3731;
  wire[46:0] T3732;
  wire[46:0] twiddle4_3_110_imag;
  wire[46:0] T3733;
  wire[46:0] T3734;
  wire[46:0] T3735;
  wire[46:0] T3736;
  wire[46:0] twiddle4_3_111_imag;
  wire[46:0] T3737;
  wire[46:0] T3738;
  wire[46:0] T3739;
  wire[46:0] T3740;
  wire T3741;
  wire T3742;
  wire T3743;
  wire T3744;
  wire[46:0] T3745;
  wire[46:0] T3746;
  wire[46:0] T3747;
  wire[46:0] T3748;
  wire[46:0] twiddle4_3_112_imag;
  wire[46:0] T3749;
  wire[46:0] T3750;
  wire[46:0] T3751;
  wire[46:0] T3752;
  wire[46:0] twiddle4_3_113_imag;
  wire[46:0] T3753;
  wire[46:0] T3754;
  wire[46:0] T3755;
  wire[46:0] T3756;
  wire T3757;
  wire[46:0] T3758;
  wire[46:0] twiddle4_3_114_imag;
  wire[46:0] T3759;
  wire[46:0] T3760;
  wire[46:0] T3761;
  wire[45:0] T3762;
  wire[45:0] T3763;
  wire T3764;
  wire[46:0] twiddle4_3_115_imag;
  wire[46:0] T3765;
  wire[46:0] T3766;
  wire[46:0] T3767;
  wire[45:0] T3768;
  wire[45:0] T3769;
  wire T3770;
  wire T3771;
  wire T3772;
  wire[46:0] T3773;
  wire[46:0] T3774;
  wire[46:0] twiddle4_3_116_imag;
  wire[46:0] T3775;
  wire[46:0] T3776;
  wire[46:0] T3777;
  wire[45:0] T3778;
  wire[45:0] T3779;
  wire T3780;
  wire[46:0] twiddle4_3_117_imag;
  wire[46:0] T3781;
  wire[46:0] T3782;
  wire[46:0] T3783;
  wire[45:0] T3784;
  wire[45:0] T3785;
  wire T3786;
  wire T3787;
  wire[46:0] T3788;
  wire[46:0] twiddle4_3_118_imag;
  wire[46:0] T3789;
  wire[46:0] T3790;
  wire[46:0] T3791;
  wire[45:0] T3792;
  wire[45:0] T3793;
  wire T3794;
  wire[46:0] twiddle4_3_119_imag;
  wire[46:0] T3795;
  wire[46:0] T3796;
  wire[46:0] T3797;
  wire[45:0] T3798;
  wire[45:0] T3799;
  wire T3800;
  wire T3801;
  wire T3802;
  wire T3803;
  wire[46:0] T3804;
  wire[46:0] T3805;
  wire[46:0] T3806;
  wire[46:0] twiddle4_3_120_imag;
  wire[46:0] T3807;
  wire[46:0] T3808;
  wire[46:0] T3809;
  wire[45:0] T3810;
  wire[45:0] T3811;
  wire T3812;
  wire[46:0] twiddle4_3_121_imag;
  wire[46:0] T3813;
  wire[46:0] T3814;
  wire[46:0] T3815;
  wire[45:0] T3816;
  wire[45:0] T3817;
  wire T3818;
  wire T3819;
  wire[46:0] T3820;
  wire[46:0] twiddle4_3_122_imag;
  wire[46:0] T3821;
  wire[46:0] T3822;
  wire[46:0] T3823;
  wire[45:0] T3824;
  wire[45:0] T3825;
  wire T3826;
  wire[46:0] twiddle4_3_123_imag;
  wire[46:0] T3827;
  wire[46:0] T3828;
  wire[46:0] T3829;
  wire[45:0] T3830;
  wire[45:0] T3831;
  wire T3832;
  wire T3833;
  wire T3834;
  wire[46:0] T3835;
  wire[46:0] T3836;
  wire[46:0] twiddle4_3_124_imag;
  wire[46:0] T3837;
  wire[46:0] T3838;
  wire[46:0] T3839;
  wire[45:0] T3840;
  wire[45:0] T3841;
  wire T3842;
  wire[46:0] twiddle4_3_125_imag;
  wire[46:0] T3843;
  wire[46:0] T3844;
  wire[46:0] T3845;
  wire[45:0] T3846;
  wire[45:0] T3847;
  wire T3848;
  wire T3849;
  wire[46:0] T3850;
  wire[46:0] twiddle4_3_126_imag;
  wire[46:0] T3851;
  wire[46:0] T3852;
  wire[46:0] T3853;
  wire[45:0] T3854;
  wire[45:0] T3855;
  wire T3856;
  wire[46:0] twiddle4_3_127_imag;
  wire[46:0] T3857;
  wire[46:0] T3858;
  wire[46:0] T3859;
  wire[45:0] T3860;
  wire[45:0] T3861;
  wire T3862;
  wire T3863;
  wire T3864;
  wire T3865;
  wire T3866;
  wire T3867;
  wire T3868;
  wire T3869;
  wire T3870;
  wire[47:0] T3871;
  wire[46:0] T3872;
  wire[46:0] T3873;
  wire[46:0] T3874;
  wire[46:0] T3875;
  wire[46:0] T3876;
  wire[46:0] T3877;
  wire[46:0] T3878;
  wire[46:0] twiddle4_3_128_imag;
  wire[46:0] T3879;
  wire[46:0] T3880;
  wire[46:0] T3881;
  wire[45:0] T3882;
  wire[45:0] T3883;
  wire T3884;
  wire[46:0] twiddle4_3_129_imag;
  wire[46:0] T3885;
  wire[46:0] T3886;
  wire[46:0] T3887;
  wire[45:0] T3888;
  wire[45:0] T3889;
  wire T3890;
  wire T3891;
  wire[46:0] T3892;
  wire[46:0] twiddle4_3_130_imag;
  wire[46:0] T3893;
  wire[46:0] T3894;
  wire[46:0] T3895;
  wire[45:0] T3896;
  wire[45:0] T3897;
  wire T3898;
  wire[46:0] twiddle4_3_131_imag;
  wire[46:0] T3899;
  wire[46:0] T3900;
  wire[46:0] T3901;
  wire[45:0] T3902;
  wire[45:0] T3903;
  wire T3904;
  wire T3905;
  wire T3906;
  wire[46:0] T3907;
  wire[46:0] T3908;
  wire[46:0] twiddle4_3_132_imag;
  wire[46:0] T3909;
  wire[46:0] T3910;
  wire[46:0] T3911;
  wire[45:0] T3912;
  wire[45:0] T3913;
  wire T3914;
  wire[46:0] twiddle4_3_133_imag;
  wire[46:0] T3915;
  wire[46:0] T3916;
  wire[46:0] T3917;
  wire[45:0] T3918;
  wire[45:0] T3919;
  wire T3920;
  wire T3921;
  wire[46:0] T3922;
  wire[46:0] twiddle4_3_134_imag;
  wire[46:0] T3923;
  wire[46:0] T3924;
  wire[46:0] T3925;
  wire[45:0] T3926;
  wire[45:0] T3927;
  wire T3928;
  wire[46:0] twiddle4_3_135_imag;
  wire[46:0] T3929;
  wire[46:0] T3930;
  wire[46:0] T3931;
  wire[45:0] T3932;
  wire[45:0] T3933;
  wire T3934;
  wire T3935;
  wire T3936;
  wire T3937;
  wire[46:0] T3938;
  wire[46:0] T3939;
  wire[46:0] T3940;
  wire[46:0] twiddle4_3_136_imag;
  wire[46:0] T3941;
  wire[46:0] T3942;
  wire[46:0] T3943;
  wire[45:0] T3944;
  wire[45:0] T3945;
  wire T3946;
  wire[46:0] twiddle4_3_137_imag;
  wire[46:0] T3947;
  wire[46:0] T3948;
  wire[46:0] T3949;
  wire[45:0] T3950;
  wire[45:0] T3951;
  wire T3952;
  wire T3953;
  wire[46:0] T3954;
  wire[46:0] twiddle4_3_138_imag;
  wire[46:0] T3955;
  wire[46:0] T3956;
  wire[46:0] T3957;
  wire[45:0] T3958;
  wire[45:0] T3959;
  wire T3960;
  wire[46:0] twiddle4_3_139_imag;
  wire[46:0] T3961;
  wire[46:0] T3962;
  wire[46:0] T3963;
  wire[45:0] T3964;
  wire[45:0] T3965;
  wire T3966;
  wire T3967;
  wire T3968;
  wire[46:0] T3969;
  wire[46:0] T3970;
  wire[46:0] twiddle4_3_140_imag;
  wire[46:0] T3971;
  wire[46:0] T3972;
  wire[46:0] T3973;
  wire[45:0] T3974;
  wire[45:0] T3975;
  wire T3976;
  wire[46:0] twiddle4_3_141_imag;
  wire[46:0] T3977;
  wire[46:0] T3978;
  wire[46:0] T3979;
  wire[45:0] T3980;
  wire[45:0] T3981;
  wire T3982;
  wire T3983;
  wire[46:0] T3984;
  wire[46:0] twiddle4_3_142_imag;
  wire[46:0] T3985;
  wire[46:0] T3986;
  wire[46:0] T3987;
  wire[45:0] T3988;
  wire[45:0] T3989;
  wire T3990;
  wire[46:0] twiddle4_3_143_imag;
  wire[46:0] T3991;
  wire[46:0] T3992;
  wire[46:0] T3993;
  wire[45:0] T3994;
  wire[45:0] T3995;
  wire T3996;
  wire T3997;
  wire T3998;
  wire T3999;
  wire T4000;
  wire[46:0] T4001;
  wire[46:0] T4002;
  wire[46:0] T4003;
  wire[46:0] T4004;
  wire[46:0] twiddle4_3_144_imag;
  wire[46:0] T4005;
  wire[46:0] T4006;
  wire[46:0] T4007;
  wire[44:0] T4008;
  wire[44:0] T4009;
  wire[1:0] T4010;
  wire T4011;
  wire[46:0] twiddle4_3_145_imag;
  wire[46:0] T4012;
  wire[46:0] T4013;
  wire[46:0] T4014;
  wire[44:0] T4015;
  wire[44:0] T4016;
  wire[1:0] T4017;
  wire T4018;
  wire T4019;
  wire[46:0] T4020;
  wire[46:0] twiddle4_3_146_imag;
  wire[46:0] T4021;
  wire[46:0] T4022;
  wire[46:0] T4023;
  wire[44:0] T4024;
  wire[44:0] T4025;
  wire[1:0] T4026;
  wire T4027;
  wire[46:0] twiddle4_3_147_imag;
  wire[46:0] T4028;
  wire[46:0] T4029;
  wire[46:0] T4030;
  wire[44:0] T4031;
  wire[44:0] T4032;
  wire[1:0] T4033;
  wire T4034;
  wire T4035;
  wire T4036;
  wire[46:0] T4037;
  wire[46:0] T4038;
  wire[46:0] twiddle4_3_148_imag;
  wire[46:0] T4039;
  wire[46:0] T4040;
  wire[46:0] T4041;
  wire[44:0] T4042;
  wire[44:0] T4043;
  wire[1:0] T4044;
  wire T4045;
  wire[46:0] twiddle4_3_149_imag;
  wire[46:0] T4046;
  wire[46:0] T4047;
  wire[46:0] T4048;
  wire[44:0] T4049;
  wire[44:0] T4050;
  wire[1:0] T4051;
  wire T4052;
  wire T4053;
  wire[46:0] T4054;
  wire[46:0] twiddle4_3_150_imag;
  wire[46:0] T4055;
  wire[46:0] T4056;
  wire[46:0] T4057;
  wire[44:0] T4058;
  wire[44:0] T4059;
  wire[1:0] T4060;
  wire T4061;
  wire[46:0] twiddle4_3_151_imag;
  wire[46:0] T4062;
  wire[46:0] T4063;
  wire[46:0] T4064;
  wire[44:0] T4065;
  wire[44:0] T4066;
  wire[1:0] T4067;
  wire T4068;
  wire T4069;
  wire T4070;
  wire T4071;
  wire[46:0] T4072;
  wire[46:0] T4073;
  wire[46:0] T4074;
  wire[46:0] twiddle4_3_152_imag;
  wire[46:0] T4075;
  wire[46:0] T4076;
  wire[46:0] T4077;
  wire[44:0] T4078;
  wire[44:0] T4079;
  wire[1:0] T4080;
  wire T4081;
  wire[46:0] twiddle4_3_153_imag;
  wire[46:0] T4082;
  wire[46:0] T4083;
  wire[46:0] T4084;
  wire[44:0] T4085;
  wire[44:0] T4086;
  wire[1:0] T4087;
  wire T4088;
  wire T4089;
  wire[46:0] T4090;
  wire[46:0] twiddle4_3_154_imag;
  wire[46:0] T4091;
  wire[46:0] T4092;
  wire[46:0] T4093;
  wire[44:0] T4094;
  wire[44:0] T4095;
  wire[1:0] T4096;
  wire T4097;
  wire[46:0] twiddle4_3_155_imag;
  wire[46:0] T4098;
  wire[46:0] T4099;
  wire[46:0] T4100;
  wire[44:0] T4101;
  wire[44:0] T4102;
  wire[1:0] T4103;
  wire T4104;
  wire T4105;
  wire T4106;
  wire[46:0] T4107;
  wire[46:0] T4108;
  wire[46:0] twiddle4_3_156_imag;
  wire[46:0] T4109;
  wire[46:0] T4110;
  wire[46:0] T4111;
  wire[44:0] T4112;
  wire[44:0] T4113;
  wire[1:0] T4114;
  wire T4115;
  wire[46:0] twiddle4_3_157_imag;
  wire[46:0] T4116;
  wire[46:0] T4117;
  wire[46:0] T4118;
  wire[44:0] T4119;
  wire[44:0] T4120;
  wire[1:0] T4121;
  wire T4122;
  wire T4123;
  wire[46:0] T4124;
  wire[46:0] twiddle4_3_158_imag;
  wire[46:0] T4125;
  wire[46:0] T4126;
  wire[46:0] T4127;
  wire[43:0] T4128;
  wire[43:0] T4129;
  wire[2:0] T4130;
  wire T4131;
  wire[46:0] twiddle4_3_159_imag;
  wire[46:0] T4132;
  wire[46:0] T4133;
  wire[46:0] T4134;
  wire[43:0] T4135;
  wire[43:0] T4136;
  wire[2:0] T4137;
  wire T4138;
  wire T4139;
  wire T4140;
  wire T4141;
  wire T4142;
  wire T4143;
  wire[46:0] T4144;
  wire[46:0] T4145;
  wire[46:0] T4146;
  wire[46:0] T4147;
  wire[46:0] T4148;
  wire[46:0] twiddle4_3_160_imag;
  wire[46:0] T4149;
  wire[46:0] T4150;
  wire[46:0] T4151;
  wire[43:0] T4152;
  wire[43:0] T4153;
  wire[2:0] T4154;
  wire T4155;
  wire[46:0] twiddle4_3_161_imag;
  wire[46:0] T4156;
  wire[46:0] T4157;
  wire[46:0] T4158;
  wire[43:0] T4159;
  wire[43:0] T4160;
  wire[2:0] T4161;
  wire T4162;
  wire T4163;
  wire[46:0] T4164;
  wire[46:0] twiddle4_3_162_imag;
  wire[46:0] T4165;
  wire[46:0] T4166;
  wire[46:0] T4167;
  wire[43:0] T4168;
  wire[43:0] T4169;
  wire[2:0] T4170;
  wire T4171;
  wire[46:0] twiddle4_3_163_imag;
  wire[46:0] T4172;
  wire[46:0] T4173;
  wire[46:0] T4174;
  wire[43:0] T4175;
  wire[43:0] T4176;
  wire[2:0] T4177;
  wire T4178;
  wire T4179;
  wire T4180;
  wire[46:0] T4181;
  wire[46:0] T4182;
  wire[46:0] twiddle4_3_164_imag;
  wire[46:0] T4183;
  wire[46:0] T4184;
  wire[46:0] T4185;
  wire[42:0] T4186;
  wire[42:0] T4187;
  wire[3:0] T4188;
  wire T4189;
  wire[46:0] twiddle4_3_165_imag;
  wire[46:0] T4190;
  wire[46:0] T4191;
  wire[46:0] T4192;
  wire[42:0] T4193;
  wire[42:0] T4194;
  wire[3:0] T4195;
  wire T4196;
  wire T4197;
  wire[46:0] T4198;
  wire[46:0] twiddle4_3_166_imag;
  wire[46:0] T4199;
  wire[46:0] T4200;
  wire[46:0] T4201;
  wire[42:0] T4202;
  wire[42:0] T4203;
  wire[3:0] T4204;
  wire T4205;
  wire[46:0] twiddle4_3_167_imag;
  wire[46:0] T4206;
  wire[46:0] T4207;
  wire[46:0] T4208;
  wire[42:0] T4209;
  wire[42:0] T4210;
  wire[3:0] T4211;
  wire T4212;
  wire T4213;
  wire T4214;
  wire T4215;
  wire[46:0] T4216;
  wire[46:0] T4217;
  wire[46:0] T4218;
  wire[46:0] twiddle4_3_168_imag;
  wire[46:0] T4219;
  wire[46:0] T4220;
  wire[46:0] T4221;
  wire[41:0] T4222;
  wire[41:0] T4223;
  wire[4:0] T4224;
  wire T4225;
  wire[46:0] twiddle4_3_169_imag;
  wire[46:0] T4226;
  wire[46:0] T4227;
  wire[46:0] T4228;
  wire[40:0] T4229;
  wire[40:0] T4230;
  wire[5:0] T4231;
  wire T4232;
  wire T4233;
  wire[46:0] T4234;
  wire[46:0] twiddle4_3_170_imag;
  wire[46:0] T4235;
  wire[46:0] T4236;
  wire[46:0] T4237;
  wire[39:0] T4238;
  wire[39:0] T4239;
  wire[6:0] T4240;
  wire T4241;
  wire[46:0] twiddle4_3_171_imag;
  wire[46:0] T4242;
  wire[46:0] T4243;
  wire[46:0] T4244;
  wire[38:0] T4245;
  wire[38:0] T4246;
  wire[7:0] T4247;
  wire T4248;
  wire T4249;
  wire T4250;
  wire[46:0] T4251;
  wire[46:0] T4252;
  wire[46:0] twiddle4_3_172_imag;
  wire[46:0] T4253;
  wire[46:0] T4254;
  wire[46:0] T4255;
  wire[40:0] T4256;
  wire[40:0] T4257;
  wire[5:0] T4258;
  wire T4259;
  wire[46:0] twiddle4_3_173_imag;
  wire[46:0] T4260;
  wire[46:0] T4261;
  wire[46:0] T4262;
  wire[41:0] T4263;
  wire[41:0] T4264;
  wire[4:0] T4265;
  wire T4266;
  wire T4267;
  wire[46:0] T4268;
  wire[46:0] twiddle4_3_174_imag;
  wire[46:0] T4269;
  wire[46:0] T4270;
  wire[46:0] T4271;
  wire[41:0] T4272;
  wire[41:0] T4273;
  wire[4:0] T4274;
  wire T4275;
  wire[46:0] twiddle4_3_175_imag;
  wire[46:0] T4276;
  wire[46:0] T4277;
  wire[46:0] T4278;
  wire[42:0] T4279;
  wire[42:0] T4280;
  wire[3:0] T4281;
  wire T4282;
  wire T4283;
  wire T4284;
  wire T4285;
  wire T4286;
  wire[46:0] T4287;
  wire[46:0] T4288;
  wire[46:0] T4289;
  wire[46:0] T4290;
  wire[46:0] twiddle4_3_176_imag;
  wire[46:0] T4291;
  wire[46:0] T4292;
  wire[46:0] T4293;
  wire[42:0] T4294;
  wire[42:0] T4295;
  wire[3:0] T4296;
  wire T4297;
  wire[46:0] twiddle4_3_177_imag;
  wire[46:0] T4298;
  wire[46:0] T4299;
  wire[46:0] T4300;
  wire[42:0] T4301;
  wire[42:0] T4302;
  wire[3:0] T4303;
  wire T4304;
  wire T4305;
  wire[46:0] T4306;
  wire[46:0] twiddle4_3_178_imag;
  wire[46:0] T4307;
  wire[46:0] T4308;
  wire[46:0] T4309;
  wire[43:0] T4310;
  wire[43:0] T4311;
  wire[2:0] T4312;
  wire T4313;
  wire[46:0] twiddle4_3_179_imag;
  wire[46:0] T4314;
  wire[46:0] T4315;
  wire[46:0] T4316;
  wire[43:0] T4317;
  wire[43:0] T4318;
  wire[2:0] T4319;
  wire T4320;
  wire T4321;
  wire T4322;
  wire[46:0] T4323;
  wire[46:0] T4324;
  wire[46:0] twiddle4_3_180_imag;
  wire[46:0] T4325;
  wire[46:0] T4326;
  wire[46:0] T4327;
  wire[43:0] T4328;
  wire[43:0] T4329;
  wire[2:0] T4330;
  wire T4331;
  wire[46:0] twiddle4_3_181_imag;
  wire[46:0] T4332;
  wire[46:0] T4333;
  wire[46:0] T4334;
  wire[43:0] T4335;
  wire[43:0] T4336;
  wire[2:0] T4337;
  wire T4338;
  wire T4339;
  wire[46:0] T4340;
  wire[46:0] twiddle4_3_182_imag;
  wire[46:0] T4341;
  wire[46:0] T4342;
  wire[46:0] T4343;
  wire[43:0] T4344;
  wire[43:0] T4345;
  wire[2:0] T4346;
  wire T4347;
  wire[46:0] twiddle4_3_183_imag;
  wire[46:0] T4348;
  wire[46:0] T4349;
  wire[46:0] T4350;
  wire[43:0] T4351;
  wire[43:0] T4352;
  wire[2:0] T4353;
  wire T4354;
  wire T4355;
  wire T4356;
  wire T4357;
  wire[46:0] T4358;
  wire[46:0] T4359;
  wire[46:0] T4360;
  wire[46:0] twiddle4_3_184_imag;
  wire[46:0] T4361;
  wire[46:0] T4362;
  wire[46:0] T4363;
  wire[43:0] T4364;
  wire[43:0] T4365;
  wire[2:0] T4366;
  wire T4367;
  wire[46:0] twiddle4_3_185_imag;
  wire[46:0] T4368;
  wire[46:0] T4369;
  wire[46:0] T4370;
  wire[44:0] T4371;
  wire[44:0] T4372;
  wire[1:0] T4373;
  wire T4374;
  wire T4375;
  wire[46:0] T4376;
  wire[46:0] twiddle4_3_186_imag;
  wire[46:0] T4377;
  wire[46:0] T4378;
  wire[46:0] T4379;
  wire[44:0] T4380;
  wire[44:0] T4381;
  wire[1:0] T4382;
  wire T4383;
  wire[46:0] twiddle4_3_187_imag;
  wire[46:0] T4384;
  wire[46:0] T4385;
  wire[46:0] T4386;
  wire[44:0] T4387;
  wire[44:0] T4388;
  wire[1:0] T4389;
  wire T4390;
  wire T4391;
  wire T4392;
  wire[46:0] T4393;
  wire[46:0] T4394;
  wire[46:0] twiddle4_3_188_imag;
  wire[46:0] T4395;
  wire[46:0] T4396;
  wire[46:0] T4397;
  wire[44:0] T4398;
  wire[44:0] T4399;
  wire[1:0] T4400;
  wire T4401;
  wire[46:0] twiddle4_3_189_imag;
  wire[46:0] T4402;
  wire[46:0] T4403;
  wire[46:0] T4404;
  wire[44:0] T4405;
  wire[44:0] T4406;
  wire[1:0] T4407;
  wire T4408;
  wire T4409;
  wire[46:0] T4410;
  wire[46:0] twiddle4_3_190_imag;
  wire[46:0] T4411;
  wire[46:0] T4412;
  wire[46:0] T4413;
  wire[44:0] T4414;
  wire[44:0] T4415;
  wire[1:0] T4416;
  wire T4417;
  wire[46:0] twiddle4_3_191_imag;
  wire[46:0] T4418;
  wire[46:0] T4419;
  wire[46:0] T4420;
  wire[44:0] T4421;
  wire[44:0] T4422;
  wire[1:0] T4423;
  wire T4424;
  wire T4425;
  wire T4426;
  wire T4427;
  wire T4428;
  wire T4429;
  wire T4430;
  wire[46:0] T4431;
  wire[46:0] T4432;
  wire[46:0] T4433;
  wire[46:0] T4434;
  wire[46:0] T4435;
  wire[46:0] T4436;
  wire[46:0] twiddle4_3_192_imag;
  wire[46:0] T4437;
  wire[46:0] T4438;
  wire[46:0] T4439;
  wire[44:0] T4440;
  wire[44:0] T4441;
  wire[1:0] T4442;
  wire T4443;
  wire[46:0] twiddle4_3_193_imag;
  wire[46:0] T4444;
  wire[46:0] T4445;
  wire[46:0] T4446;
  wire[44:0] T4447;
  wire[44:0] T4448;
  wire[1:0] T4449;
  wire T4450;
  wire T4451;
  wire[46:0] T4452;
  wire[46:0] twiddle4_3_194_imag;
  wire[46:0] T4453;
  wire[46:0] T4454;
  wire[46:0] T4455;
  wire[44:0] T4456;
  wire[44:0] T4457;
  wire[1:0] T4458;
  wire T4459;
  wire[46:0] twiddle4_3_195_imag;
  wire[46:0] T4460;
  wire[46:0] T4461;
  wire[46:0] T4462;
  wire[44:0] T4463;
  wire[44:0] T4464;
  wire[1:0] T4465;
  wire T4466;
  wire T4467;
  wire T4468;
  wire[46:0] T4469;
  wire[46:0] T4470;
  wire[46:0] twiddle4_3_196_imag;
  wire[46:0] T4471;
  wire[46:0] T4472;
  wire[46:0] T4473;
  wire[44:0] T4474;
  wire[44:0] T4475;
  wire[1:0] T4476;
  wire T4477;
  wire[46:0] twiddle4_3_197_imag;
  wire[46:0] T4478;
  wire[46:0] T4479;
  wire[46:0] T4480;
  wire[44:0] T4481;
  wire[44:0] T4482;
  wire[1:0] T4483;
  wire T4484;
  wire T4485;
  wire[46:0] T4486;
  wire[46:0] twiddle4_3_198_imag;
  wire[46:0] T4487;
  wire[46:0] T4488;
  wire[46:0] T4489;
  wire[44:0] T4490;
  wire[44:0] T4491;
  wire[1:0] T4492;
  wire T4493;
  wire[46:0] twiddle4_3_199_imag;
  wire[46:0] T4494;
  wire[46:0] T4495;
  wire[46:0] T4496;
  wire[45:0] T4497;
  wire[45:0] T4498;
  wire T4499;
  wire T4500;
  wire T4501;
  wire T4502;
  wire[46:0] T4503;
  wire[46:0] T4504;
  wire[46:0] T4505;
  wire[46:0] twiddle4_3_200_imag;
  wire[46:0] T4506;
  wire[46:0] T4507;
  wire[46:0] T4508;
  wire[45:0] T4509;
  wire[45:0] T4510;
  wire T4511;
  wire[46:0] twiddle4_3_201_imag;
  wire[46:0] T4512;
  wire[46:0] T4513;
  wire[46:0] T4514;
  wire[45:0] T4515;
  wire[45:0] T4516;
  wire T4517;
  wire T4518;
  wire[46:0] T4519;
  wire[46:0] twiddle4_3_202_imag;
  wire[46:0] T4520;
  wire[46:0] T4521;
  wire[46:0] T4522;
  wire[45:0] T4523;
  wire[45:0] T4524;
  wire T4525;
  wire[46:0] twiddle4_3_203_imag;
  wire[46:0] T4526;
  wire[46:0] T4527;
  wire[46:0] T4528;
  wire[45:0] T4529;
  wire[45:0] T4530;
  wire T4531;
  wire T4532;
  wire T4533;
  wire[46:0] T4534;
  wire[46:0] T4535;
  wire[46:0] twiddle4_3_204_imag;
  wire[46:0] T4536;
  wire[46:0] T4537;
  wire[46:0] T4538;
  wire[45:0] T4539;
  wire[45:0] T4540;
  wire T4541;
  wire[46:0] twiddle4_3_205_imag;
  wire[46:0] T4542;
  wire[46:0] T4543;
  wire[46:0] T4544;
  wire[45:0] T4545;
  wire[45:0] T4546;
  wire T4547;
  wire T4548;
  wire[46:0] T4549;
  wire[46:0] twiddle4_3_206_imag;
  wire[46:0] T4550;
  wire[46:0] T4551;
  wire[46:0] T4552;
  wire[45:0] T4553;
  wire[45:0] T4554;
  wire T4555;
  wire[46:0] twiddle4_3_207_imag;
  wire[46:0] T4556;
  wire[46:0] T4557;
  wire[46:0] T4558;
  wire[45:0] T4559;
  wire[45:0] T4560;
  wire T4561;
  wire T4562;
  wire T4563;
  wire T4564;
  wire T4565;
  wire[46:0] T4566;
  wire[46:0] T4567;
  wire[46:0] T4568;
  wire[46:0] T4569;
  wire[46:0] twiddle4_3_208_imag;
  wire[46:0] T4570;
  wire[46:0] T4571;
  wire[46:0] T4572;
  wire[45:0] T4573;
  wire[45:0] T4574;
  wire T4575;
  wire[46:0] twiddle4_3_209_imag;
  wire[46:0] T4576;
  wire[46:0] T4577;
  wire[46:0] T4578;
  wire[45:0] T4579;
  wire[45:0] T4580;
  wire T4581;
  wire T4582;
  wire[46:0] T4583;
  wire[46:0] twiddle4_3_210_imag;
  wire[46:0] T4584;
  wire[46:0] T4585;
  wire[46:0] T4586;
  wire[45:0] T4587;
  wire[45:0] T4588;
  wire T4589;
  wire[46:0] twiddle4_3_211_imag;
  wire[46:0] T4590;
  wire[46:0] T4591;
  wire[46:0] T4592;
  wire[45:0] T4593;
  wire[45:0] T4594;
  wire T4595;
  wire T4596;
  wire T4597;
  wire[46:0] T4598;
  wire[46:0] T4599;
  wire[46:0] twiddle4_3_212_imag;
  wire[46:0] T4600;
  wire[46:0] T4601;
  wire[46:0] T4602;
  wire[45:0] T4603;
  wire[45:0] T4604;
  wire T4605;
  wire[46:0] twiddle4_3_213_imag;
  wire[46:0] T4606;
  wire[46:0] T4607;
  wire[46:0] T4608;
  wire[45:0] T4609;
  wire[45:0] T4610;
  wire T4611;
  wire T4612;
  wire[46:0] T4613;
  wire[46:0] twiddle4_3_214_imag;
  wire[46:0] T4614;
  wire[46:0] T4615;
  wire[46:0] T4616;
  wire[45:0] T4617;
  wire[45:0] T4618;
  wire T4619;
  wire[46:0] twiddle4_3_215_imag;
  wire[46:0] T4620;
  wire[46:0] T4621;
  wire[46:0] T4622;
  wire[45:0] T4623;
  wire[45:0] T4624;
  wire T4625;
  wire T4626;
  wire T4627;
  wire T4628;
  wire[46:0] T4629;
  wire[46:0] T4630;
  wire[46:0] T4631;
  wire[46:0] twiddle4_3_216_imag;
  wire[46:0] T4632;
  wire[46:0] T4633;
  wire[46:0] T4634;
  wire[45:0] T4635;
  wire[45:0] T4636;
  wire T4637;
  wire[46:0] twiddle4_3_217_imag;
  wire[46:0] T4638;
  wire[46:0] T4639;
  wire[46:0] T4640;
  wire[45:0] T4641;
  wire[45:0] T4642;
  wire T4643;
  wire T4644;
  wire[46:0] T4645;
  wire[46:0] twiddle4_3_218_imag;
  wire[46:0] T4646;
  wire[46:0] T4647;
  wire[46:0] T4648;
  wire[45:0] T4649;
  wire[45:0] T4650;
  wire T4651;
  wire[46:0] twiddle4_3_219_imag;
  wire[46:0] T4652;
  wire[46:0] T4653;
  wire[46:0] T4654;
  wire[45:0] T4655;
  wire[45:0] T4656;
  wire T4657;
  wire T4658;
  wire T4659;
  wire[46:0] T4660;
  wire[46:0] T4661;
  wire[46:0] twiddle4_3_220_imag;
  wire[46:0] T4662;
  wire[46:0] T4663;
  wire[46:0] T4664;
  wire[45:0] T4665;
  wire[45:0] T4666;
  wire T4667;
  wire[46:0] twiddle4_3_221_imag;
  wire[46:0] T4668;
  wire[46:0] T4669;
  wire[46:0] T4670;
  wire[45:0] T4671;
  wire[45:0] T4672;
  wire T4673;
  wire T4674;
  wire[46:0] T4675;
  wire[46:0] twiddle4_3_222_imag;
  wire[46:0] T4676;
  wire[46:0] T4677;
  wire[46:0] T4678;
  wire[45:0] T4679;
  wire[45:0] T4680;
  wire T4681;
  wire[46:0] twiddle4_3_223_imag;
  wire[46:0] T4682;
  wire[46:0] T4683;
  wire[46:0] T4684;
  wire[45:0] T4685;
  wire[45:0] T4686;
  wire T4687;
  wire T4688;
  wire T4689;
  wire T4690;
  wire T4691;
  wire T4692;
  wire[46:0] T4693;
  wire[46:0] T4694;
  wire[46:0] T4695;
  wire[46:0] T4696;
  wire[46:0] T4697;
  wire[46:0] twiddle4_3_224_imag;
  wire[46:0] T4698;
  wire[46:0] T4699;
  wire[46:0] T4700;
  wire[45:0] T4701;
  wire[45:0] T4702;
  wire T4703;
  wire[46:0] twiddle4_3_225_imag;
  wire[46:0] T4704;
  wire[46:0] T4705;
  wire[46:0] T4706;
  wire[45:0] T4707;
  wire[45:0] T4708;
  wire T4709;
  wire T4710;
  wire[46:0] T4711;
  wire[46:0] twiddle4_3_226_imag;
  wire[46:0] T4712;
  wire[46:0] T4713;
  wire[46:0] T4714;
  wire[45:0] T4715;
  wire[45:0] T4716;
  wire T4717;
  wire[46:0] twiddle4_3_227_imag;
  wire[46:0] T4718;
  wire[46:0] T4719;
  wire[46:0] T4720;
  wire[45:0] T4721;
  wire[45:0] T4722;
  wire T4723;
  wire T4724;
  wire T4725;
  wire[46:0] T4726;
  wire[46:0] T4727;
  wire[46:0] twiddle4_3_228_imag;
  wire[46:0] T4728;
  wire[46:0] T4729;
  wire[46:0] T4730;
  wire[46:0] T4731;
  wire[46:0] twiddle4_3_229_imag;
  wire[46:0] T4732;
  wire[46:0] T4733;
  wire[46:0] T4734;
  wire[46:0] T4735;
  wire T4736;
  wire[46:0] T4737;
  wire[46:0] twiddle4_3_230_imag;
  wire[46:0] T4738;
  wire[46:0] T4739;
  wire[46:0] T4740;
  wire[46:0] T4741;
  wire[46:0] twiddle4_3_231_imag;
  wire[46:0] T4742;
  wire[46:0] T4743;
  wire[46:0] T4744;
  wire[46:0] T4745;
  wire T4746;
  wire T4747;
  wire T4748;
  wire[46:0] T4749;
  wire[46:0] T4750;
  wire[46:0] T4751;
  wire[46:0] twiddle4_3_232_imag;
  wire[46:0] T4752;
  wire[46:0] T4753;
  wire[46:0] T4754;
  wire[46:0] T4755;
  wire[46:0] twiddle4_3_233_imag;
  wire[46:0] T4756;
  wire[46:0] T4757;
  wire[46:0] T4758;
  wire[46:0] T4759;
  wire T4760;
  wire[46:0] T4761;
  wire[46:0] twiddle4_3_234_imag;
  wire[46:0] T4762;
  wire[46:0] T4763;
  wire[46:0] T4764;
  wire[46:0] T4765;
  wire[46:0] twiddle4_3_235_imag;
  wire[46:0] T4766;
  wire[46:0] T4767;
  wire[46:0] T4768;
  wire[46:0] T4769;
  wire T4770;
  wire T4771;
  wire[46:0] T4772;
  wire[46:0] T4773;
  wire[46:0] twiddle4_3_236_imag;
  wire[46:0] T4774;
  wire[46:0] T4775;
  wire[46:0] T4776;
  wire[46:0] T4777;
  wire[46:0] twiddle4_3_237_imag;
  wire[46:0] T4778;
  wire[46:0] T4779;
  wire[46:0] T4780;
  wire[46:0] T4781;
  wire T4782;
  wire[46:0] T4783;
  wire[46:0] twiddle4_3_238_imag;
  wire[46:0] T4784;
  wire[46:0] T4785;
  wire[46:0] T4786;
  wire[46:0] T4787;
  wire[46:0] twiddle4_3_239_imag;
  wire[46:0] T4788;
  wire[46:0] T4789;
  wire[46:0] T4790;
  wire[46:0] T4791;
  wire T4792;
  wire T4793;
  wire T4794;
  wire T4795;
  wire[46:0] T4796;
  wire[46:0] T4797;
  wire[46:0] T4798;
  wire[46:0] T4799;
  wire[46:0] twiddle4_3_240_imag;
  wire[46:0] T4800;
  wire[46:0] T4801;
  wire[46:0] T4802;
  wire[46:0] T4803;
  wire[46:0] twiddle4_3_241_imag;
  wire[46:0] T4804;
  wire[46:0] T4805;
  wire[46:0] T4806;
  wire[46:0] T4807;
  wire T4808;
  wire[46:0] T4809;
  wire[46:0] twiddle4_3_242_imag;
  wire[46:0] T4810;
  wire[46:0] T4811;
  wire[46:0] T4812;
  wire[46:0] T4813;
  wire[46:0] twiddle4_3_243_imag;
  wire[46:0] T4814;
  wire[46:0] T4815;
  wire[46:0] T4816;
  wire[46:0] T4817;
  wire T4818;
  wire T4819;
  wire[46:0] T4820;
  wire[46:0] T4821;
  wire[46:0] twiddle4_3_244_imag;
  wire[46:0] T4822;
  wire[46:0] T4823;
  wire[46:0] T4824;
  wire[46:0] T4825;
  wire[46:0] twiddle4_3_245_imag;
  wire[46:0] T4826;
  wire[46:0] T4827;
  wire[46:0] T4828;
  wire[46:0] T4829;
  wire T4830;
  wire[46:0] T4831;
  wire[46:0] twiddle4_3_246_imag;
  wire[46:0] T4832;
  wire[46:0] T4833;
  wire[46:0] T4834;
  wire[46:0] T4835;
  wire[46:0] twiddle4_3_247_imag;
  wire[46:0] T4836;
  wire[46:0] T4837;
  wire[46:0] T4838;
  wire[46:0] T4839;
  wire T4840;
  wire T4841;
  wire T4842;
  wire[46:0] T4843;
  wire[46:0] T4844;
  wire[46:0] T4845;
  wire[46:0] twiddle4_3_248_imag;
  wire[46:0] T4846;
  wire[46:0] T4847;
  wire[46:0] T4848;
  wire[46:0] T4849;
  wire[46:0] twiddle4_3_249_imag;
  wire[46:0] T4850;
  wire[46:0] T4851;
  wire[46:0] T4852;
  wire[46:0] T4853;
  wire T4854;
  wire[46:0] T4855;
  wire[46:0] twiddle4_3_250_imag;
  wire[46:0] T4856;
  wire[46:0] T4857;
  wire[46:0] T4858;
  wire[46:0] T4859;
  wire[46:0] twiddle4_3_251_imag;
  wire[46:0] T4860;
  wire[46:0] T4861;
  wire[46:0] T4862;
  wire[46:0] T4863;
  wire T4864;
  wire T4865;
  wire[46:0] T4866;
  wire[46:0] T4867;
  wire[46:0] twiddle4_3_252_imag;
  wire[46:0] T4868;
  wire[46:0] T4869;
  wire[46:0] T4870;
  wire[46:0] T4871;
  wire[46:0] twiddle4_3_253_imag;
  wire[46:0] T4872;
  wire[46:0] T4873;
  wire[46:0] T4874;
  wire[46:0] T4875;
  wire T4876;
  wire[46:0] T4877;
  wire[46:0] twiddle4_3_254_imag;
  wire[46:0] T4878;
  wire[46:0] T4879;
  wire[46:0] T4880;
  wire[46:0] T4881;
  wire[46:0] twiddle4_3_255_imag;
  wire[46:0] T4882;
  wire[46:0] T4883;
  wire[46:0] T4884;
  wire[46:0] T4885;
  wire T4886;
  wire T4887;
  wire T4888;
  wire T4889;
  wire T4890;
  wire T4891;
  wire T4892;
  wire T4893;
  wire T4894;
  wire[47:0] T4895;
  wire[46:0] T4896;
  wire[46:0] T4897;
  wire[46:0] T4898;
  wire[46:0] T4899;
  wire[46:0] T4900;
  wire[46:0] T4901;
  wire[46:0] T4902;
  wire[46:0] T4903;
  wire[46:0] twiddle4_3_256_imag;
  wire[46:0] T4904;
  wire[46:0] T4905;
  wire[46:0] T4906;
  wire[46:0] T4907;
  wire[46:0] twiddle4_3_257_imag;
  wire[46:0] T4908;
  wire[46:0] T4909;
  wire[46:0] T4910;
  wire[46:0] T4911;
  wire T4912;
  wire[46:0] T4913;
  wire[46:0] twiddle4_3_258_imag;
  wire[46:0] T4914;
  wire[46:0] T4915;
  wire[46:0] T4916;
  wire[46:0] T4917;
  wire[46:0] twiddle4_3_259_imag;
  wire[46:0] T4918;
  wire[46:0] T4919;
  wire[46:0] T4920;
  wire[46:0] T4921;
  wire T4922;
  wire T4923;
  wire[46:0] T4924;
  wire[46:0] T4925;
  wire[46:0] twiddle4_3_260_imag;
  wire[46:0] T4926;
  wire[46:0] T4927;
  wire[46:0] T4928;
  wire[46:0] T4929;
  wire[46:0] twiddle4_3_261_imag;
  wire[46:0] T4930;
  wire[46:0] T4931;
  wire[46:0] T4932;
  wire[46:0] T4933;
  wire T4934;
  wire[46:0] T4935;
  wire[46:0] twiddle4_3_262_imag;
  wire[46:0] T4936;
  wire[46:0] T4937;
  wire[46:0] T4938;
  wire[46:0] T4939;
  wire[46:0] twiddle4_3_263_imag;
  wire[46:0] T4940;
  wire[46:0] T4941;
  wire[46:0] T4942;
  wire[46:0] T4943;
  wire T4944;
  wire T4945;
  wire T4946;
  wire[46:0] T4947;
  wire[46:0] T4948;
  wire[46:0] T4949;
  wire[46:0] twiddle4_3_264_imag;
  wire[46:0] T4950;
  wire[46:0] T4951;
  wire[46:0] T4952;
  wire[46:0] T4953;
  wire[46:0] twiddle4_3_265_imag;
  wire[46:0] T4954;
  wire[46:0] T4955;
  wire[46:0] T4956;
  wire[46:0] T4957;
  wire T4958;
  wire[46:0] T4959;
  wire[46:0] twiddle4_3_266_imag;
  wire[46:0] T4960;
  wire[46:0] T4961;
  wire[46:0] T4962;
  wire[46:0] T4963;
  wire[46:0] twiddle4_3_267_imag;
  wire[46:0] T4964;
  wire[46:0] T4965;
  wire[46:0] T4966;
  wire[46:0] T4967;
  wire T4968;
  wire T4969;
  wire[46:0] T4970;
  wire[46:0] T4971;
  wire[46:0] twiddle4_3_268_imag;
  wire[46:0] T4972;
  wire[46:0] T4973;
  wire[46:0] T4974;
  wire[46:0] T4975;
  wire[46:0] twiddle4_3_269_imag;
  wire[46:0] T4976;
  wire[46:0] T4977;
  wire[46:0] T4978;
  wire[46:0] T4979;
  wire T4980;
  wire[46:0] T4981;
  wire[46:0] twiddle4_3_270_imag;
  wire[46:0] T4982;
  wire[46:0] T4983;
  wire[46:0] T4984;
  wire[46:0] T4985;
  wire[46:0] twiddle4_3_271_imag;
  wire[46:0] T4986;
  wire[46:0] T4987;
  wire[46:0] T4988;
  wire[46:0] T4989;
  wire T4990;
  wire T4991;
  wire T4992;
  wire T4993;
  wire[46:0] T4994;
  wire[46:0] T4995;
  wire[46:0] T4996;
  wire[46:0] T4997;
  wire[46:0] twiddle4_3_272_imag;
  wire[46:0] T4998;
  wire[46:0] T4999;
  wire[46:0] T5000;
  wire[46:0] T5001;
  wire[46:0] twiddle4_3_273_imag;
  wire[46:0] T5002;
  wire[46:0] T5003;
  wire[46:0] T5004;
  wire[46:0] T5005;
  wire T5006;
  wire[46:0] T5007;
  wire[46:0] twiddle4_3_274_imag;
  wire[46:0] T5008;
  wire[46:0] T5009;
  wire[46:0] T5010;
  wire[46:0] T5011;
  wire[46:0] twiddle4_3_275_imag;
  wire[46:0] T5012;
  wire[46:0] T5013;
  wire[46:0] T5014;
  wire[46:0] T5015;
  wire T5016;
  wire T5017;
  wire[46:0] T5018;
  wire[46:0] T5019;
  wire[46:0] twiddle4_3_276_imag;
  wire[46:0] T5020;
  wire[46:0] T5021;
  wire[46:0] T5022;
  wire[46:0] T5023;
  wire[46:0] twiddle4_3_277_imag;
  wire[46:0] T5024;
  wire[46:0] T5025;
  wire[46:0] T5026;
  wire[46:0] T5027;
  wire T5028;
  wire[46:0] T5029;
  wire[46:0] twiddle4_3_278_imag;
  wire[46:0] T5030;
  wire[46:0] T5031;
  wire[46:0] T5032;
  wire[46:0] T5033;
  wire[46:0] twiddle4_3_279_imag;
  wire[46:0] T5034;
  wire[46:0] T5035;
  wire[46:0] T5036;
  wire[46:0] T5037;
  wire T5038;
  wire T5039;
  wire T5040;
  wire[46:0] T5041;
  wire[46:0] T5042;
  wire[46:0] T5043;
  wire[46:0] twiddle4_3_280_imag;
  wire[46:0] T5044;
  wire[46:0] T5045;
  wire[46:0] T5046;
  wire[46:0] T5047;
  wire[46:0] twiddle4_3_281_imag;
  wire[46:0] T5048;
  wire[46:0] T5049;
  wire[46:0] T5050;
  wire[46:0] T5051;
  wire T5052;
  wire[46:0] T5053;
  wire[46:0] twiddle4_3_282_imag;
  wire[46:0] T5054;
  wire[46:0] T5055;
  wire[46:0] T5056;
  wire[46:0] T5057;
  wire[46:0] twiddle4_3_283_imag;
  wire[46:0] T5058;
  wire[46:0] T5059;
  wire[46:0] T5060;
  wire[46:0] T5061;
  wire T5062;
  wire T5063;
  wire[46:0] T5064;
  wire[46:0] T5065;
  wire[46:0] twiddle4_3_284_imag;
  wire[46:0] T5066;
  wire[46:0] T5067;
  wire[46:0] T5068;
  wire[46:0] T5069;
  wire[46:0] twiddle4_3_285_imag;
  wire[46:0] T5070;
  wire[45:0] T5071;
  wire[45:0] T5072;
  wire T5073;
  wire[46:0] T5074;
  wire[46:0] T5075;
  wire T5076;
  wire[46:0] T5077;
  wire[46:0] twiddle4_3_286_imag;
  wire[46:0] T5078;
  wire[45:0] T5079;
  wire[45:0] T5080;
  wire T5081;
  wire[46:0] T5082;
  wire[46:0] T5083;
  wire[46:0] twiddle4_3_287_imag;
  wire[46:0] T5084;
  wire[45:0] T5085;
  wire[45:0] T5086;
  wire T5087;
  wire[46:0] T5088;
  wire[46:0] T5089;
  wire T5090;
  wire T5091;
  wire T5092;
  wire T5093;
  wire T5094;
  wire[46:0] T5095;
  wire[46:0] T5096;
  wire[46:0] T5097;
  wire[46:0] T5098;
  wire[46:0] T5099;
  wire[46:0] twiddle4_3_288_imag;
  wire[46:0] T5100;
  wire[45:0] T5101;
  wire[45:0] T5102;
  wire T5103;
  wire[46:0] T5104;
  wire[46:0] T5105;
  wire[46:0] twiddle4_3_289_imag;
  wire[46:0] T5106;
  wire[45:0] T5107;
  wire[45:0] T5108;
  wire T5109;
  wire[46:0] T5110;
  wire[46:0] T5111;
  wire T5112;
  wire[46:0] T5113;
  wire[46:0] twiddle4_3_290_imag;
  wire[46:0] T5114;
  wire[45:0] T5115;
  wire[45:0] T5116;
  wire T5117;
  wire[46:0] T5118;
  wire[46:0] T5119;
  wire[46:0] twiddle4_3_291_imag;
  wire[46:0] T5120;
  wire[45:0] T5121;
  wire[45:0] T5122;
  wire T5123;
  wire[46:0] T5124;
  wire[46:0] T5125;
  wire T5126;
  wire T5127;
  wire[46:0] T5128;
  wire[46:0] T5129;
  wire[46:0] twiddle4_3_292_imag;
  wire[46:0] T5130;
  wire[45:0] T5131;
  wire[45:0] T5132;
  wire T5133;
  wire[46:0] T5134;
  wire[46:0] T5135;
  wire[46:0] twiddle4_3_293_imag;
  wire[46:0] T5136;
  wire[45:0] T5137;
  wire[45:0] T5138;
  wire T5139;
  wire[46:0] T5140;
  wire[46:0] T5141;
  wire T5142;
  wire[46:0] T5143;
  wire[46:0] twiddle4_3_294_imag;
  wire[46:0] T5144;
  wire[45:0] T5145;
  wire[45:0] T5146;
  wire T5147;
  wire[46:0] T5148;
  wire[46:0] T5149;
  wire[46:0] twiddle4_3_295_imag;
  wire[46:0] T5150;
  wire[45:0] T5151;
  wire[45:0] T5152;
  wire T5153;
  wire[46:0] T5154;
  wire[46:0] T5155;
  wire T5156;
  wire T5157;
  wire T5158;
  wire[46:0] T5159;
  wire[46:0] T5160;
  wire[46:0] T5161;
  wire[46:0] twiddle4_3_296_imag;
  wire[46:0] T5162;
  wire[45:0] T5163;
  wire[45:0] T5164;
  wire T5165;
  wire[46:0] T5166;
  wire[46:0] T5167;
  wire[46:0] twiddle4_3_297_imag;
  wire[46:0] T5168;
  wire[45:0] T5169;
  wire[45:0] T5170;
  wire T5171;
  wire[46:0] T5172;
  wire[46:0] T5173;
  wire T5174;
  wire[46:0] T5175;
  wire[46:0] twiddle4_3_298_imag;
  wire[46:0] T5176;
  wire[45:0] T5177;
  wire[45:0] T5178;
  wire T5179;
  wire[46:0] T5180;
  wire[46:0] T5181;
  wire[46:0] twiddle4_3_299_imag;
  wire[46:0] T5182;
  wire[45:0] T5183;
  wire[45:0] T5184;
  wire T5185;
  wire[46:0] T5186;
  wire[46:0] T5187;
  wire T5188;
  wire T5189;
  wire[46:0] T5190;
  wire[46:0] T5191;
  wire[46:0] twiddle4_3_300_imag;
  wire[46:0] T5192;
  wire[45:0] T5193;
  wire[45:0] T5194;
  wire T5195;
  wire[46:0] T5196;
  wire[46:0] T5197;
  wire[46:0] twiddle4_3_301_imag;
  wire[46:0] T5198;
  wire[45:0] T5199;
  wire[45:0] T5200;
  wire T5201;
  wire[46:0] T5202;
  wire[46:0] T5203;
  wire T5204;
  wire[46:0] T5205;
  wire[46:0] twiddle4_3_302_imag;
  wire[46:0] T5206;
  wire[45:0] T5207;
  wire[45:0] T5208;
  wire T5209;
  wire[46:0] T5210;
  wire[46:0] T5211;
  wire[46:0] twiddle4_3_303_imag;
  wire[46:0] T5212;
  wire[45:0] T5213;
  wire[45:0] T5214;
  wire T5215;
  wire[46:0] T5216;
  wire[46:0] T5217;
  wire T5218;
  wire T5219;
  wire T5220;
  wire T5221;
  wire[46:0] T5222;
  wire[46:0] T5223;
  wire[46:0] T5224;
  wire[46:0] T5225;
  wire[46:0] twiddle4_3_304_imag;
  wire[46:0] T5226;
  wire[45:0] T5227;
  wire[45:0] T5228;
  wire T5229;
  wire[46:0] T5230;
  wire[46:0] T5231;
  wire[46:0] twiddle4_3_305_imag;
  wire[46:0] T5232;
  wire[45:0] T5233;
  wire[45:0] T5234;
  wire T5235;
  wire[46:0] T5236;
  wire[46:0] T5237;
  wire T5238;
  wire[46:0] T5239;
  wire[46:0] twiddle4_3_306_imag;
  wire[46:0] T5240;
  wire[45:0] T5241;
  wire[45:0] T5242;
  wire T5243;
  wire[46:0] T5244;
  wire[46:0] T5245;
  wire[46:0] twiddle4_3_307_imag;
  wire[46:0] T5246;
  wire[45:0] T5247;
  wire[45:0] T5248;
  wire T5249;
  wire[46:0] T5250;
  wire[46:0] T5251;
  wire T5252;
  wire T5253;
  wire[46:0] T5254;
  wire[46:0] T5255;
  wire[46:0] twiddle4_3_308_imag;
  wire[46:0] T5256;
  wire[45:0] T5257;
  wire[45:0] T5258;
  wire T5259;
  wire[46:0] T5260;
  wire[46:0] T5261;
  wire[46:0] twiddle4_3_309_imag;
  wire[46:0] T5262;
  wire[45:0] T5263;
  wire[45:0] T5264;
  wire T5265;
  wire[46:0] T5266;
  wire[46:0] T5267;
  wire T5268;
  wire[46:0] T5269;
  wire[46:0] twiddle4_3_310_imag;
  wire[46:0] T5270;
  wire[45:0] T5271;
  wire[45:0] T5272;
  wire T5273;
  wire[46:0] T5274;
  wire[46:0] T5275;
  wire[46:0] twiddle4_3_311_imag;
  wire[46:0] T5276;
  wire[45:0] T5277;
  wire[45:0] T5278;
  wire T5279;
  wire[46:0] T5280;
  wire[46:0] T5281;
  wire T5282;
  wire T5283;
  wire T5284;
  wire[46:0] T5285;
  wire[46:0] T5286;
  wire[46:0] T5287;
  wire[46:0] twiddle4_3_312_imag;
  wire[46:0] T5288;
  wire[45:0] T5289;
  wire[45:0] T5290;
  wire T5291;
  wire[46:0] T5292;
  wire[46:0] T5293;
  wire[46:0] twiddle4_3_313_imag;
  wire[46:0] T5294;
  wire[45:0] T5295;
  wire[45:0] T5296;
  wire T5297;
  wire[46:0] T5298;
  wire[46:0] T5299;
  wire T5300;
  wire[46:0] T5301;
  wire[46:0] twiddle4_3_314_imag;
  wire[46:0] T5302;
  wire[44:0] T5303;
  wire[44:0] T5304;
  wire[1:0] T5305;
  wire T5306;
  wire[46:0] T5307;
  wire[46:0] T5308;
  wire[46:0] twiddle4_3_315_imag;
  wire[46:0] T5309;
  wire[44:0] T5310;
  wire[44:0] T5311;
  wire[1:0] T5312;
  wire T5313;
  wire[46:0] T5314;
  wire[46:0] T5315;
  wire T5316;
  wire T5317;
  wire[46:0] T5318;
  wire[46:0] T5319;
  wire[46:0] twiddle4_3_316_imag;
  wire[46:0] T5320;
  wire[44:0] T5321;
  wire[44:0] T5322;
  wire[1:0] T5323;
  wire T5324;
  wire[46:0] T5325;
  wire[46:0] T5326;
  wire[46:0] twiddle4_3_317_imag;
  wire[46:0] T5327;
  wire[44:0] T5328;
  wire[44:0] T5329;
  wire[1:0] T5330;
  wire T5331;
  wire[46:0] T5332;
  wire[46:0] T5333;
  wire T5334;
  wire[46:0] T5335;
  wire[46:0] twiddle4_3_318_imag;
  wire[46:0] T5336;
  wire[44:0] T5337;
  wire[44:0] T5338;
  wire[1:0] T5339;
  wire T5340;
  wire[46:0] T5341;
  wire[46:0] T5342;
  wire[46:0] twiddle4_3_319_imag;
  wire[46:0] T5343;
  wire[44:0] T5344;
  wire[44:0] T5345;
  wire[1:0] T5346;
  wire T5347;
  wire[46:0] T5348;
  wire[46:0] T5349;
  wire T5350;
  wire T5351;
  wire T5352;
  wire T5353;
  wire T5354;
  wire T5355;
  wire[46:0] T5356;
  wire[46:0] T5357;
  wire[46:0] T5358;
  wire[46:0] T5359;
  wire[46:0] T5360;
  wire[46:0] T5361;
  wire[46:0] twiddle4_3_320_imag;
  wire[46:0] T5362;
  wire[44:0] T5363;
  wire[44:0] T5364;
  wire[1:0] T5365;
  wire T5366;
  wire[46:0] T5367;
  wire[46:0] T5368;
  wire[46:0] twiddle4_3_321_imag;
  wire[46:0] T5369;
  wire[44:0] T5370;
  wire[44:0] T5371;
  wire[1:0] T5372;
  wire T5373;
  wire[46:0] T5374;
  wire[46:0] T5375;
  wire T5376;
  wire[46:0] T5377;
  wire[46:0] twiddle4_3_322_imag;
  wire[46:0] T5378;
  wire[44:0] T5379;
  wire[44:0] T5380;
  wire[1:0] T5381;
  wire T5382;
  wire[46:0] T5383;
  wire[46:0] T5384;
  wire[46:0] twiddle4_3_323_imag;
  wire[46:0] T5385;
  wire[44:0] T5386;
  wire[44:0] T5387;
  wire[1:0] T5388;
  wire T5389;
  wire[46:0] T5390;
  wire[46:0] T5391;
  wire T5392;
  wire T5393;
  wire[46:0] T5394;
  wire[46:0] T5395;
  wire[46:0] twiddle4_3_324_imag;
  wire[46:0] T5396;
  wire[44:0] T5397;
  wire[44:0] T5398;
  wire[1:0] T5399;
  wire T5400;
  wire[46:0] T5401;
  wire[46:0] T5402;
  wire[46:0] twiddle4_3_325_imag;
  wire[46:0] T5403;
  wire[44:0] T5404;
  wire[44:0] T5405;
  wire[1:0] T5406;
  wire T5407;
  wire[46:0] T5408;
  wire[46:0] T5409;
  wire T5410;
  wire[46:0] T5411;
  wire[46:0] twiddle4_3_326_imag;
  wire[46:0] T5412;
  wire[44:0] T5413;
  wire[44:0] T5414;
  wire[1:0] T5415;
  wire T5416;
  wire[46:0] T5417;
  wire[46:0] T5418;
  wire[46:0] twiddle4_3_327_imag;
  wire[46:0] T5419;
  wire[44:0] T5420;
  wire[44:0] T5421;
  wire[1:0] T5422;
  wire T5423;
  wire[46:0] T5424;
  wire[46:0] T5425;
  wire T5426;
  wire T5427;
  wire T5428;
  wire[46:0] T5429;
  wire[46:0] T5430;
  wire[46:0] T5431;
  wire[46:0] twiddle4_3_328_imag;
  wire[46:0] T5432;
  wire[43:0] T5433;
  wire[43:0] T5434;
  wire[2:0] T5435;
  wire T5436;
  wire[46:0] T5437;
  wire[46:0] T5438;
  wire[46:0] twiddle4_3_329_imag;
  wire[46:0] T5439;
  wire[43:0] T5440;
  wire[43:0] T5441;
  wire[2:0] T5442;
  wire T5443;
  wire[46:0] T5444;
  wire[46:0] T5445;
  wire T5446;
  wire[46:0] T5447;
  wire[46:0] twiddle4_3_330_imag;
  wire[46:0] T5448;
  wire[43:0] T5449;
  wire[43:0] T5450;
  wire[2:0] T5451;
  wire T5452;
  wire[46:0] T5453;
  wire[46:0] T5454;
  wire[46:0] twiddle4_3_331_imag;
  wire[46:0] T5455;
  wire[43:0] T5456;
  wire[43:0] T5457;
  wire[2:0] T5458;
  wire T5459;
  wire[46:0] T5460;
  wire[46:0] T5461;
  wire T5462;
  wire T5463;
  wire[46:0] T5464;
  wire[46:0] T5465;
  wire[46:0] twiddle4_3_332_imag;
  wire[46:0] T5466;
  wire[43:0] T5467;
  wire[43:0] T5468;
  wire[2:0] T5469;
  wire T5470;
  wire[46:0] T5471;
  wire[46:0] T5472;
  wire[46:0] twiddle4_3_333_imag;
  wire[46:0] T5473;
  wire[43:0] T5474;
  wire[43:0] T5475;
  wire[2:0] T5476;
  wire T5477;
  wire[46:0] T5478;
  wire[46:0] T5479;
  wire T5480;
  wire[46:0] T5481;
  wire[46:0] twiddle4_3_334_imag;
  wire[46:0] T5482;
  wire[43:0] T5483;
  wire[43:0] T5484;
  wire[2:0] T5485;
  wire T5486;
  wire[46:0] T5487;
  wire[46:0] T5488;
  wire[46:0] twiddle4_3_335_imag;
  wire[46:0] T5489;
  wire[42:0] T5490;
  wire[42:0] T5491;
  wire[3:0] T5492;
  wire T5493;
  wire[46:0] T5494;
  wire[46:0] T5495;
  wire T5496;
  wire T5497;
  wire T5498;
  wire T5499;
  wire[46:0] T5500;
  wire[46:0] T5501;
  wire[46:0] T5502;
  wire[46:0] T5503;
  wire[46:0] twiddle4_3_336_imag;
  wire[46:0] T5504;
  wire[42:0] T5505;
  wire[42:0] T5506;
  wire[3:0] T5507;
  wire T5508;
  wire[46:0] T5509;
  wire[46:0] T5510;
  wire[46:0] twiddle4_3_337_imag;
  wire[46:0] T5511;
  wire[42:0] T5512;
  wire[42:0] T5513;
  wire[3:0] T5514;
  wire T5515;
  wire[46:0] T5516;
  wire[46:0] T5517;
  wire T5518;
  wire[46:0] T5519;
  wire[46:0] twiddle4_3_338_imag;
  wire[46:0] T5520;
  wire[41:0] T5521;
  wire[41:0] T5522;
  wire[4:0] T5523;
  wire T5524;
  wire[46:0] T5525;
  wire[46:0] T5526;
  wire[46:0] twiddle4_3_339_imag;
  wire[46:0] T5527;
  wire[41:0] T5528;
  wire[41:0] T5529;
  wire[4:0] T5530;
  wire T5531;
  wire[46:0] T5532;
  wire[46:0] T5533;
  wire T5534;
  wire T5535;
  wire[46:0] T5536;
  wire[46:0] T5537;
  wire[46:0] twiddle4_3_340_imag;
  wire[46:0] T5538;
  wire[40:0] T5539;
  wire[40:0] T5540;
  wire[5:0] T5541;
  wire T5542;
  wire[46:0] T5543;
  wire[46:0] T5544;
  wire[46:0] twiddle4_3_341_imag;
  wire[46:0] T5545;
  wire[38:0] T5546;
  wire[38:0] T5547;
  wire[7:0] T5548;
  wire T5549;
  wire[46:0] T5550;
  wire[46:0] T5551;
  wire T5552;
  wire[46:0] T5553;
  wire[46:0] twiddle4_3_342_imag;
  wire[46:0] T5554;
  wire[39:0] T5555;
  wire[39:0] T5556;
  wire[6:0] T5557;
  wire T5558;
  wire[46:0] T5559;
  wire[46:0] T5560;
  wire[46:0] twiddle4_3_343_imag;
  wire[46:0] T5561;
  wire[40:0] T5562;
  wire[40:0] T5563;
  wire[5:0] T5564;
  wire T5565;
  wire[46:0] T5566;
  wire[46:0] T5567;
  wire T5568;
  wire T5569;
  wire T5570;
  wire[46:0] T5571;
  wire[46:0] T5572;
  wire[46:0] T5573;
  wire[46:0] twiddle4_3_344_imag;
  wire[46:0] T5574;
  wire[41:0] T5575;
  wire[41:0] T5576;
  wire[4:0] T5577;
  wire T5578;
  wire[46:0] T5579;
  wire[46:0] T5580;
  wire[46:0] twiddle4_3_345_imag;
  wire[46:0] T5581;
  wire[42:0] T5582;
  wire[42:0] T5583;
  wire[3:0] T5584;
  wire T5585;
  wire[46:0] T5586;
  wire[46:0] T5587;
  wire T5588;
  wire[46:0] T5589;
  wire[46:0] twiddle4_3_346_imag;
  wire[46:0] T5590;
  wire[42:0] T5591;
  wire[42:0] T5592;
  wire[3:0] T5593;
  wire T5594;
  wire[46:0] T5595;
  wire[46:0] T5596;
  wire[46:0] twiddle4_3_347_imag;
  wire[46:0] T5597;
  wire[42:0] T5598;
  wire[42:0] T5599;
  wire[3:0] T5600;
  wire T5601;
  wire[46:0] T5602;
  wire[46:0] T5603;
  wire T5604;
  wire T5605;
  wire[46:0] T5606;
  wire[46:0] T5607;
  wire[46:0] twiddle4_3_348_imag;
  wire[46:0] T5608;
  wire[42:0] T5609;
  wire[42:0] T5610;
  wire[3:0] T5611;
  wire T5612;
  wire[46:0] T5613;
  wire[46:0] T5614;
  wire[46:0] twiddle4_3_349_imag;
  wire[46:0] T5615;
  wire[43:0] T5616;
  wire[43:0] T5617;
  wire[2:0] T5618;
  wire T5619;
  wire[46:0] T5620;
  wire[46:0] T5621;
  wire T5622;
  wire[46:0] T5623;
  wire[46:0] twiddle4_3_350_imag;
  wire[46:0] T5624;
  wire[43:0] T5625;
  wire[43:0] T5626;
  wire[2:0] T5627;
  wire T5628;
  wire[46:0] T5629;
  wire[46:0] T5630;
  wire[46:0] twiddle4_3_351_imag;
  wire[46:0] T5631;
  wire[43:0] T5632;
  wire[43:0] T5633;
  wire[2:0] T5634;
  wire T5635;
  wire[46:0] T5636;
  wire[46:0] T5637;
  wire T5638;
  wire T5639;
  wire T5640;
  wire T5641;
  wire T5642;
  wire[46:0] T5643;
  wire[46:0] T5644;
  wire[46:0] T5645;
  wire[46:0] T5646;
  wire[46:0] T5647;
  wire[46:0] twiddle4_3_352_imag;
  wire[46:0] T5648;
  wire[43:0] T5649;
  wire[43:0] T5650;
  wire[2:0] T5651;
  wire T5652;
  wire[46:0] T5653;
  wire[46:0] T5654;
  wire[46:0] twiddle4_3_353_imag;
  wire[46:0] T5655;
  wire[43:0] T5656;
  wire[43:0] T5657;
  wire[2:0] T5658;
  wire T5659;
  wire[46:0] T5660;
  wire[46:0] T5661;
  wire T5662;
  wire[46:0] T5663;
  wire[46:0] twiddle4_3_354_imag;
  wire[46:0] T5664;
  wire[43:0] T5665;
  wire[43:0] T5666;
  wire[2:0] T5667;
  wire T5668;
  wire[46:0] T5669;
  wire[46:0] T5670;
  wire[46:0] twiddle4_3_355_imag;
  wire[46:0] T5671;
  wire[44:0] T5672;
  wire[44:0] T5673;
  wire[1:0] T5674;
  wire T5675;
  wire[46:0] T5676;
  wire[46:0] T5677;
  wire T5678;
  wire T5679;
  wire[46:0] T5680;
  wire[46:0] T5681;
  wire[46:0] twiddle4_3_356_imag;
  wire[46:0] T5682;
  wire[44:0] T5683;
  wire[44:0] T5684;
  wire[1:0] T5685;
  wire T5686;
  wire[46:0] T5687;
  wire[46:0] T5688;
  wire[46:0] twiddle4_3_357_imag;
  wire[46:0] T5689;
  wire[44:0] T5690;
  wire[44:0] T5691;
  wire[1:0] T5692;
  wire T5693;
  wire[46:0] T5694;
  wire[46:0] T5695;
  wire T5696;
  wire[46:0] T5697;
  wire[46:0] twiddle4_3_358_imag;
  wire[46:0] T5698;
  wire[44:0] T5699;
  wire[44:0] T5700;
  wire[1:0] T5701;
  wire T5702;
  wire[46:0] T5703;
  wire[46:0] T5704;
  wire[46:0] twiddle4_3_359_imag;
  wire[46:0] T5705;
  wire[44:0] T5706;
  wire[44:0] T5707;
  wire[1:0] T5708;
  wire T5709;
  wire[46:0] T5710;
  wire[46:0] T5711;
  wire T5712;
  wire T5713;
  wire T5714;
  wire[46:0] T5715;
  wire[46:0] T5716;
  wire[46:0] T5717;
  wire[46:0] twiddle4_3_360_imag;
  wire[46:0] T5718;
  wire[44:0] T5719;
  wire[44:0] T5720;
  wire[1:0] T5721;
  wire T5722;
  wire[46:0] T5723;
  wire[46:0] T5724;
  wire[46:0] twiddle4_3_361_imag;
  wire[46:0] T5725;
  wire[44:0] T5726;
  wire[44:0] T5727;
  wire[1:0] T5728;
  wire T5729;
  wire[46:0] T5730;
  wire[46:0] T5731;
  wire T5732;
  wire[46:0] T5733;
  wire[46:0] twiddle4_3_362_imag;
  wire[46:0] T5734;
  wire[44:0] T5735;
  wire[44:0] T5736;
  wire[1:0] T5737;
  wire T5738;
  wire[46:0] T5739;
  wire[46:0] T5740;
  wire[46:0] twiddle4_3_363_imag;
  wire[46:0] T5741;
  wire[44:0] T5742;
  wire[44:0] T5743;
  wire[1:0] T5744;
  wire T5745;
  wire[46:0] T5746;
  wire[46:0] T5747;
  wire T5748;
  wire T5749;
  wire[46:0] T5750;
  wire[46:0] T5751;
  wire[46:0] twiddle4_3_364_imag;
  wire[46:0] T5752;
  wire[44:0] T5753;
  wire[44:0] T5754;
  wire[1:0] T5755;
  wire T5756;
  wire[46:0] T5757;
  wire[46:0] T5758;
  wire[46:0] twiddle4_3_365_imag;
  wire[46:0] T5759;
  wire[44:0] T5760;
  wire[44:0] T5761;
  wire[1:0] T5762;
  wire T5763;
  wire[46:0] T5764;
  wire[46:0] T5765;
  wire T5766;
  wire[46:0] T5767;
  wire[46:0] twiddle4_3_366_imag;
  wire[46:0] T5768;
  wire[44:0] T5769;
  wire[44:0] T5770;
  wire[1:0] T5771;
  wire T5772;
  wire[46:0] T5773;
  wire[46:0] T5774;
  wire[46:0] twiddle4_3_367_imag;
  wire[46:0] T5775;
  wire[44:0] T5776;
  wire[44:0] T5777;
  wire[1:0] T5778;
  wire T5779;
  wire[46:0] T5780;
  wire[46:0] T5781;
  wire T5782;
  wire T5783;
  wire T5784;
  wire T5785;
  wire[46:0] T5786;
  wire[46:0] T5787;
  wire[46:0] T5788;
  wire[46:0] T5789;
  wire[46:0] twiddle4_3_368_imag;
  wire[46:0] T5790;
  wire[44:0] T5791;
  wire[44:0] T5792;
  wire[1:0] T5793;
  wire T5794;
  wire[46:0] T5795;
  wire[46:0] T5796;
  wire[46:0] twiddle4_3_369_imag;
  wire[46:0] T5797;
  wire[45:0] T5798;
  wire[45:0] T5799;
  wire T5800;
  wire[46:0] T5801;
  wire[46:0] T5802;
  wire T5803;
  wire[46:0] T5804;
  wire[46:0] twiddle4_3_370_imag;
  wire[46:0] T5805;
  wire[45:0] T5806;
  wire[45:0] T5807;
  wire T5808;
  wire[46:0] T5809;
  wire[46:0] T5810;
  wire[46:0] twiddle4_3_371_imag;
  wire[46:0] T5811;
  wire[45:0] T5812;
  wire[45:0] T5813;
  wire T5814;
  wire[46:0] T5815;
  wire[46:0] T5816;
  wire T5817;
  wire T5818;
  wire[46:0] T5819;
  wire[46:0] T5820;
  wire[46:0] twiddle4_3_372_imag;
  wire[46:0] T5821;
  wire[45:0] T5822;
  wire[45:0] T5823;
  wire T5824;
  wire[46:0] T5825;
  wire[46:0] T5826;
  wire[46:0] twiddle4_3_373_imag;
  wire[46:0] T5827;
  wire[45:0] T5828;
  wire[45:0] T5829;
  wire T5830;
  wire[46:0] T5831;
  wire[46:0] T5832;
  wire T5833;
  wire[46:0] T5834;
  wire[46:0] twiddle4_3_374_imag;
  wire[46:0] T5835;
  wire[45:0] T5836;
  wire[45:0] T5837;
  wire T5838;
  wire[46:0] T5839;
  wire[46:0] T5840;
  wire[46:0] twiddle4_3_375_imag;
  wire[46:0] T5841;
  wire[45:0] T5842;
  wire[45:0] T5843;
  wire T5844;
  wire[46:0] T5845;
  wire[46:0] T5846;
  wire T5847;
  wire T5848;
  wire T5849;
  wire[46:0] T5850;
  wire[46:0] T5851;
  wire[46:0] T5852;
  wire[46:0] twiddle4_3_376_imag;
  wire[46:0] T5853;
  wire[45:0] T5854;
  wire[45:0] T5855;
  wire T5856;
  wire[46:0] T5857;
  wire[46:0] T5858;
  wire[46:0] twiddle4_3_377_imag;
  wire[46:0] T5859;
  wire[45:0] T5860;
  wire[45:0] T5861;
  wire T5862;
  wire[46:0] T5863;
  wire[46:0] T5864;
  wire T5865;
  wire[46:0] T5866;
  wire[46:0] twiddle4_3_378_imag;
  wire[46:0] T5867;
  wire[45:0] T5868;
  wire[45:0] T5869;
  wire T5870;
  wire[46:0] T5871;
  wire[46:0] T5872;
  wire[46:0] twiddle4_3_379_imag;
  wire[46:0] T5873;
  wire[45:0] T5874;
  wire[45:0] T5875;
  wire T5876;
  wire[46:0] T5877;
  wire[46:0] T5878;
  wire T5879;
  wire T5880;
  wire[46:0] T5881;
  wire[46:0] T5882;
  wire[46:0] twiddle4_3_380_imag;
  wire[46:0] T5883;
  wire[45:0] T5884;
  wire[45:0] T5885;
  wire T5886;
  wire[46:0] T5887;
  wire[46:0] T5888;
  wire[46:0] twiddle4_3_381_imag;
  wire[46:0] T5889;
  wire[45:0] T5890;
  wire[45:0] T5891;
  wire T5892;
  wire[46:0] T5893;
  wire[46:0] T5894;
  wire T5895;
  wire[46:0] T5896;
  wire[46:0] twiddle4_3_382_imag;
  wire[46:0] T5897;
  wire[45:0] T5898;
  wire[45:0] T5899;
  wire T5900;
  wire[46:0] T5901;
  wire[46:0] T5902;
  wire[46:0] twiddle4_3_383_imag;
  wire[46:0] T5903;
  wire[45:0] T5904;
  wire[45:0] T5905;
  wire T5906;
  wire[46:0] T5907;
  wire[46:0] T5908;
  wire T5909;
  wire T5910;
  wire T5911;
  wire T5912;
  wire T5913;
  wire T5914;
  wire T5915;
  wire[46:0] T5916;
  wire[46:0] T5917;
  wire[46:0] T5918;
  wire[46:0] T5919;
  wire[46:0] T5920;
  wire[46:0] T5921;
  wire[46:0] T5922;
  wire[46:0] twiddle4_3_384_imag;
  wire[46:0] T5923;
  wire[45:0] T5924;
  wire[45:0] T5925;
  wire T5926;
  wire[46:0] T5927;
  wire[46:0] T5928;
  wire[46:0] twiddle4_3_385_imag;
  wire[46:0] T5929;
  wire[45:0] T5930;
  wire[45:0] T5931;
  wire T5932;
  wire[46:0] T5933;
  wire[46:0] T5934;
  wire T5935;
  wire[46:0] T5936;
  wire[46:0] twiddle4_3_386_imag;
  wire[46:0] T5937;
  wire[45:0] T5938;
  wire[45:0] T5939;
  wire T5940;
  wire[46:0] T5941;
  wire[46:0] T5942;
  wire[46:0] twiddle4_3_387_imag;
  wire[46:0] T5943;
  wire[45:0] T5944;
  wire[45:0] T5945;
  wire T5946;
  wire[46:0] T5947;
  wire[46:0] T5948;
  wire T5949;
  wire T5950;
  wire[46:0] T5951;
  wire[46:0] T5952;
  wire[46:0] twiddle4_3_388_imag;
  wire[46:0] T5953;
  wire[45:0] T5954;
  wire[45:0] T5955;
  wire T5956;
  wire[46:0] T5957;
  wire[46:0] T5958;
  wire[46:0] twiddle4_3_389_imag;
  wire[46:0] T5959;
  wire[45:0] T5960;
  wire[45:0] T5961;
  wire T5962;
  wire[46:0] T5963;
  wire[46:0] T5964;
  wire T5965;
  wire[46:0] T5966;
  wire[46:0] twiddle4_3_390_imag;
  wire[46:0] T5967;
  wire[45:0] T5968;
  wire[45:0] T5969;
  wire T5970;
  wire[46:0] T5971;
  wire[46:0] T5972;
  wire[46:0] twiddle4_3_391_imag;
  wire[46:0] T5973;
  wire[45:0] T5974;
  wire[45:0] T5975;
  wire T5976;
  wire[46:0] T5977;
  wire[46:0] T5978;
  wire T5979;
  wire T5980;
  wire T5981;
  wire[46:0] T5982;
  wire[46:0] T5983;
  wire[46:0] T5984;
  wire[46:0] twiddle4_3_392_imag;
  wire[46:0] T5985;
  wire[45:0] T5986;
  wire[45:0] T5987;
  wire T5988;
  wire[46:0] T5989;
  wire[46:0] T5990;
  wire[46:0] twiddle4_3_393_imag;
  wire[46:0] T5991;
  wire[45:0] T5992;
  wire[45:0] T5993;
  wire T5994;
  wire[46:0] T5995;
  wire[46:0] T5996;
  wire T5997;
  wire[46:0] T5998;
  wire[46:0] twiddle4_3_394_imag;
  wire[46:0] T5999;
  wire[45:0] T6000;
  wire[45:0] T6001;
  wire T6002;
  wire[46:0] T6003;
  wire[46:0] T6004;
  wire[46:0] twiddle4_3_395_imag;
  wire[46:0] T6005;
  wire[45:0] T6006;
  wire[45:0] T6007;
  wire T6008;
  wire[46:0] T6009;
  wire[46:0] T6010;
  wire T6011;
  wire T6012;
  wire[46:0] T6013;
  wire[46:0] T6014;
  wire[46:0] twiddle4_3_396_imag;
  wire[46:0] T6015;
  wire[45:0] T6016;
  wire[45:0] T6017;
  wire T6018;
  wire[46:0] T6019;
  wire[46:0] T6020;
  wire[46:0] twiddle4_3_397_imag;
  wire[46:0] T6021;
  wire[45:0] T6022;
  wire[45:0] T6023;
  wire T6024;
  wire[46:0] T6025;
  wire[46:0] T6026;
  wire T6027;
  wire[46:0] T6028;
  wire[46:0] twiddle4_3_398_imag;
  wire[46:0] T6029;
  wire[45:0] T6030;
  wire[45:0] T6031;
  wire T6032;
  wire[46:0] T6033;
  wire[46:0] T6034;
  wire[46:0] twiddle4_3_399_imag;
  wire[46:0] T6035;
  wire[46:0] T6036;
  wire[46:0] T6037;
  wire[46:0] T6038;
  wire T6039;
  wire T6040;
  wire T6041;
  wire T6042;
  wire[46:0] T6043;
  wire[46:0] T6044;
  wire[46:0] T6045;
  wire[46:0] T6046;
  wire[46:0] twiddle4_3_400_imag;
  wire[46:0] T6047;
  wire[46:0] T6048;
  wire[46:0] T6049;
  wire[46:0] T6050;
  wire[46:0] twiddle4_3_401_imag;
  wire[46:0] T6051;
  wire[46:0] T6052;
  wire[46:0] T6053;
  wire[46:0] T6054;
  wire T6055;
  wire[46:0] T6056;
  wire[46:0] twiddle4_3_402_imag;
  wire[46:0] T6057;
  wire[46:0] T6058;
  wire[46:0] T6059;
  wire[46:0] T6060;
  wire[46:0] twiddle4_3_403_imag;
  wire[46:0] T6061;
  wire[46:0] T6062;
  wire[46:0] T6063;
  wire[46:0] T6064;
  wire T6065;
  wire T6066;
  wire[46:0] T6067;
  wire[46:0] T6068;
  wire[46:0] twiddle4_3_404_imag;
  wire[46:0] T6069;
  wire[46:0] T6070;
  wire[46:0] T6071;
  wire[46:0] T6072;
  wire[46:0] twiddle4_3_405_imag;
  wire[46:0] T6073;
  wire[46:0] T6074;
  wire[46:0] T6075;
  wire[46:0] T6076;
  wire T6077;
  wire[46:0] T6078;
  wire[46:0] twiddle4_3_406_imag;
  wire[46:0] T6079;
  wire[46:0] T6080;
  wire[46:0] T6081;
  wire[46:0] T6082;
  wire[46:0] twiddle4_3_407_imag;
  wire[46:0] T6083;
  wire[46:0] T6084;
  wire[46:0] T6085;
  wire[46:0] T6086;
  wire T6087;
  wire T6088;
  wire T6089;
  wire[46:0] T6090;
  wire[46:0] T6091;
  wire[46:0] T6092;
  wire[46:0] twiddle4_3_408_imag;
  wire[46:0] T6093;
  wire[46:0] T6094;
  wire[46:0] T6095;
  wire[46:0] T6096;
  wire[46:0] twiddle4_3_409_imag;
  wire[46:0] T6097;
  wire[46:0] T6098;
  wire[46:0] T6099;
  wire[46:0] T6100;
  wire T6101;
  wire[46:0] T6102;
  wire[46:0] twiddle4_3_410_imag;
  wire[46:0] T6103;
  wire[46:0] T6104;
  wire[46:0] T6105;
  wire[46:0] T6106;
  wire[46:0] twiddle4_3_411_imag;
  wire[46:0] T6107;
  wire[46:0] T6108;
  wire[46:0] T6109;
  wire[46:0] T6110;
  wire T6111;
  wire T6112;
  wire[46:0] T6113;
  wire[46:0] T6114;
  wire[46:0] twiddle4_3_412_imag;
  wire[46:0] T6115;
  wire[46:0] T6116;
  wire[46:0] T6117;
  wire[46:0] T6118;
  wire[46:0] twiddle4_3_413_imag;
  wire[46:0] T6119;
  wire[46:0] T6120;
  wire[46:0] T6121;
  wire[46:0] T6122;
  wire T6123;
  wire[46:0] T6124;
  wire[46:0] twiddle4_3_414_imag;
  wire[46:0] T6125;
  wire[46:0] T6126;
  wire[46:0] T6127;
  wire[46:0] T6128;
  wire[46:0] twiddle4_3_415_imag;
  wire[46:0] T6129;
  wire[46:0] T6130;
  wire[46:0] T6131;
  wire[46:0] T6132;
  wire T6133;
  wire T6134;
  wire T6135;
  wire T6136;
  wire T6137;
  wire[46:0] T6138;
  wire[46:0] T6139;
  wire[46:0] T6140;
  wire[46:0] T6141;
  wire[46:0] T6142;
  wire[46:0] twiddle4_3_416_imag;
  wire[46:0] T6143;
  wire[46:0] T6144;
  wire[46:0] T6145;
  wire[46:0] T6146;
  wire[46:0] twiddle4_3_417_imag;
  wire[46:0] T6147;
  wire[46:0] T6148;
  wire[46:0] T6149;
  wire[46:0] T6150;
  wire T6151;
  wire[46:0] T6152;
  wire[46:0] twiddle4_3_418_imag;
  wire[46:0] T6153;
  wire[46:0] T6154;
  wire[46:0] T6155;
  wire[46:0] T6156;
  wire[46:0] twiddle4_3_419_imag;
  wire[46:0] T6157;
  wire[46:0] T6158;
  wire[46:0] T6159;
  wire[46:0] T6160;
  wire T6161;
  wire T6162;
  wire[46:0] T6163;
  wire[46:0] T6164;
  wire[46:0] twiddle4_3_420_imag;
  wire[46:0] T6165;
  wire[46:0] T6166;
  wire[46:0] T6167;
  wire[46:0] T6168;
  wire[46:0] twiddle4_3_421_imag;
  wire[46:0] T6169;
  wire[46:0] T6170;
  wire[46:0] T6171;
  wire[46:0] T6172;
  wire T6173;
  wire[46:0] T6174;
  wire[46:0] twiddle4_3_422_imag;
  wire[46:0] T6175;
  wire[46:0] T6176;
  wire[46:0] T6177;
  wire[46:0] T6178;
  wire[46:0] twiddle4_3_423_imag;
  wire[46:0] T6179;
  wire[46:0] T6180;
  wire[46:0] T6181;
  wire[46:0] T6182;
  wire T6183;
  wire T6184;
  wire T6185;
  wire[46:0] T6186;
  wire[46:0] T6187;
  wire[46:0] T6188;
  wire[46:0] twiddle4_3_424_imag;
  wire[46:0] T6189;
  wire[46:0] T6190;
  wire[46:0] T6191;
  wire[46:0] T6192;
  wire[46:0] twiddle4_3_425_imag;
  wire[46:0] T6193;
  wire[46:0] T6194;
  wire[46:0] T6195;
  wire[46:0] T6196;
  wire T6197;
  wire[46:0] T6198;
  wire[46:0] twiddle4_3_426_imag;
  wire[46:0] T6199;
  wire[46:0] T6200;
  wire[46:0] T6201;
  wire[46:0] T6202;
  wire[46:0] twiddle4_3_427_imag;
  wire[46:0] T6203;
  wire[46:0] T6204;
  wire[46:0] T6205;
  wire[46:0] T6206;
  wire T6207;
  wire T6208;
  wire[46:0] T6209;
  wire[46:0] T6210;
  wire[46:0] twiddle4_3_428_imag;
  wire[46:0] T6211;
  wire[46:0] T6212;
  wire[46:0] T6213;
  wire[46:0] T6214;
  wire[46:0] twiddle4_3_429_imag;
  wire[46:0] T6215;
  wire[46:0] T6216;
  wire[46:0] T6217;
  wire[46:0] T6218;
  wire T6219;
  wire[46:0] T6220;
  wire[46:0] twiddle4_3_430_imag;
  wire[46:0] T6221;
  wire[46:0] T6222;
  wire[46:0] T6223;
  wire[46:0] T6224;
  wire[46:0] twiddle4_3_431_imag;
  wire[46:0] T6225;
  wire[46:0] T6226;
  wire[46:0] T6227;
  wire[46:0] T6228;
  wire T6229;
  wire T6230;
  wire T6231;
  wire T6232;
  wire[46:0] T6233;
  wire[46:0] T6234;
  wire[46:0] T6235;
  wire[46:0] T6236;
  wire[46:0] twiddle4_3_432_imag;
  wire[46:0] T6237;
  wire[46:0] T6238;
  wire[46:0] T6239;
  wire[46:0] T6240;
  wire[46:0] twiddle4_3_433_imag;
  wire[46:0] T6241;
  wire[46:0] T6242;
  wire[46:0] T6243;
  wire[46:0] T6244;
  wire T6245;
  wire[46:0] T6246;
  wire[46:0] twiddle4_3_434_imag;
  wire[46:0] T6247;
  wire[46:0] T6248;
  wire[46:0] T6249;
  wire[46:0] T6250;
  wire[46:0] twiddle4_3_435_imag;
  wire[46:0] T6251;
  wire[46:0] T6252;
  wire[46:0] T6253;
  wire[46:0] T6254;
  wire T6255;
  wire T6256;
  wire[46:0] T6257;
  wire[46:0] T6258;
  wire[46:0] twiddle4_3_436_imag;
  wire[46:0] T6259;
  wire[46:0] T6260;
  wire[46:0] T6261;
  wire[46:0] T6262;
  wire[46:0] twiddle4_3_437_imag;
  wire[46:0] T6263;
  wire[46:0] T6264;
  wire[46:0] T6265;
  wire[46:0] T6266;
  wire T6267;
  wire[46:0] T6268;
  wire[46:0] twiddle4_3_438_imag;
  wire[46:0] T6269;
  wire[46:0] T6270;
  wire[46:0] T6271;
  wire[46:0] T6272;
  wire[46:0] twiddle4_3_439_imag;
  wire[46:0] T6273;
  wire[46:0] T6274;
  wire[46:0] T6275;
  wire[46:0] T6276;
  wire T6277;
  wire T6278;
  wire T6279;
  wire[46:0] T6280;
  wire[46:0] T6281;
  wire[46:0] T6282;
  wire[46:0] twiddle4_3_440_imag;
  wire[46:0] T6283;
  wire[46:0] T6284;
  wire[46:0] T6285;
  wire[46:0] T6286;
  wire[46:0] twiddle4_3_441_imag;
  wire[46:0] T6287;
  wire[46:0] T6288;
  wire[46:0] T6289;
  wire[46:0] T6290;
  wire T6291;
  wire[46:0] T6292;
  wire[46:0] twiddle4_3_442_imag;
  wire[46:0] T6293;
  wire[46:0] T6294;
  wire[46:0] T6295;
  wire[46:0] T6296;
  wire[46:0] twiddle4_3_443_imag;
  wire[46:0] T6297;
  wire[46:0] T6298;
  wire[46:0] T6299;
  wire[46:0] T6300;
  wire T6301;
  wire T6302;
  wire[46:0] T6303;
  wire[46:0] T6304;
  wire[46:0] twiddle4_3_444_imag;
  wire[46:0] T6305;
  wire[46:0] T6306;
  wire[46:0] T6307;
  wire[46:0] T6308;
  wire[46:0] twiddle4_3_445_imag;
  wire[46:0] T6309;
  wire[46:0] T6310;
  wire[46:0] T6311;
  wire[46:0] T6312;
  wire T6313;
  wire[46:0] T6314;
  wire[46:0] twiddle4_3_446_imag;
  wire[46:0] T6315;
  wire[46:0] T6316;
  wire[46:0] T6317;
  wire[46:0] T6318;
  wire[46:0] twiddle4_3_447_imag;
  wire[46:0] T6319;
  wire[46:0] T6320;
  wire[46:0] T6321;
  wire[46:0] T6322;
  wire T6323;
  wire T6324;
  wire T6325;
  wire T6326;
  wire T6327;
  wire T6328;
  wire[46:0] T6329;
  wire[46:0] T6330;
  wire[46:0] T6331;
  wire[46:0] T6332;
  wire[46:0] T6333;
  wire[46:0] T6334;
  wire[46:0] twiddle4_3_448_imag;
  wire[46:0] T6335;
  wire[46:0] T6336;
  wire[46:0] T6337;
  wire[46:0] T6338;
  wire[46:0] twiddle4_3_449_imag;
  wire[46:0] T6339;
  wire[46:0] T6340;
  wire[46:0] T6341;
  wire[46:0] T6342;
  wire T6343;
  wire[46:0] T6344;
  wire[46:0] twiddle4_3_450_imag;
  wire[46:0] T6345;
  wire[46:0] T6346;
  wire[46:0] T6347;
  wire[46:0] T6348;
  wire[46:0] twiddle4_3_451_imag;
  wire[46:0] T6349;
  wire[46:0] T6350;
  wire[46:0] T6351;
  wire[46:0] T6352;
  wire T6353;
  wire T6354;
  wire[46:0] T6355;
  wire[46:0] T6356;
  wire[46:0] twiddle4_3_452_imag;
  wire[46:0] T6357;
  wire[46:0] T6358;
  wire[46:0] T6359;
  wire[46:0] T6360;
  wire[46:0] twiddle4_3_453_imag;
  wire[46:0] T6361;
  wire[46:0] T6362;
  wire[46:0] T6363;
  wire[46:0] T6364;
  wire T6365;
  wire[46:0] T6366;
  wire[46:0] twiddle4_3_454_imag;
  wire[46:0] T6367;
  wire[46:0] T6368;
  wire[46:0] T6369;
  wire[46:0] T6370;
  wire[46:0] twiddle4_3_455_imag;
  wire[46:0] T6371;
  wire[46:0] T6372;
  wire[46:0] T6373;
  wire[46:0] T6374;
  wire T6375;
  wire T6376;
  wire T6377;
  wire[46:0] T6378;
  wire[46:0] T6379;
  wire[46:0] T6380;
  wire[46:0] twiddle4_3_456_imag;
  wire[46:0] T6381;
  wire[46:0] T6382;
  wire[46:0] T6383;
  wire[45:0] T6384;
  wire[45:0] T6385;
  wire T6386;
  wire[46:0] twiddle4_3_457_imag;
  wire[46:0] T6387;
  wire[46:0] T6388;
  wire[46:0] T6389;
  wire[45:0] T6390;
  wire[45:0] T6391;
  wire T6392;
  wire T6393;
  wire[46:0] T6394;
  wire[46:0] twiddle4_3_458_imag;
  wire[46:0] T6395;
  wire[46:0] T6396;
  wire[46:0] T6397;
  wire[45:0] T6398;
  wire[45:0] T6399;
  wire T6400;
  wire[46:0] twiddle4_3_459_imag;
  wire[46:0] T6401;
  wire[46:0] T6402;
  wire[46:0] T6403;
  wire[45:0] T6404;
  wire[45:0] T6405;
  wire T6406;
  wire T6407;
  wire T6408;
  wire[46:0] T6409;
  wire[46:0] T6410;
  wire[46:0] twiddle4_3_460_imag;
  wire[46:0] T6411;
  wire[46:0] T6412;
  wire[46:0] T6413;
  wire[45:0] T6414;
  wire[45:0] T6415;
  wire T6416;
  wire[46:0] twiddle4_3_461_imag;
  wire[46:0] T6417;
  wire[46:0] T6418;
  wire[46:0] T6419;
  wire[45:0] T6420;
  wire[45:0] T6421;
  wire T6422;
  wire T6423;
  wire[46:0] T6424;
  wire[46:0] twiddle4_3_462_imag;
  wire[46:0] T6425;
  wire[46:0] T6426;
  wire[46:0] T6427;
  wire[45:0] T6428;
  wire[45:0] T6429;
  wire T6430;
  wire[46:0] twiddle4_3_463_imag;
  wire[46:0] T6431;
  wire[46:0] T6432;
  wire[46:0] T6433;
  wire[45:0] T6434;
  wire[45:0] T6435;
  wire T6436;
  wire T6437;
  wire T6438;
  wire T6439;
  wire T6440;
  wire[46:0] T6441;
  wire[46:0] T6442;
  wire[46:0] T6443;
  wire[46:0] T6444;
  wire[46:0] twiddle4_3_464_imag;
  wire[46:0] T6445;
  wire[46:0] T6446;
  wire[46:0] T6447;
  wire[45:0] T6448;
  wire[45:0] T6449;
  wire T6450;
  wire[46:0] twiddle4_3_465_imag;
  wire[46:0] T6451;
  wire[46:0] T6452;
  wire[46:0] T6453;
  wire[45:0] T6454;
  wire[45:0] T6455;
  wire T6456;
  wire T6457;
  wire[46:0] T6458;
  wire[46:0] twiddle4_3_466_imag;
  wire[46:0] T6459;
  wire[46:0] T6460;
  wire[46:0] T6461;
  wire[45:0] T6462;
  wire[45:0] T6463;
  wire T6464;
  wire[46:0] twiddle4_3_467_imag;
  wire[46:0] T6465;
  wire[46:0] T6466;
  wire[46:0] T6467;
  wire[45:0] T6468;
  wire[45:0] T6469;
  wire T6470;
  wire T6471;
  wire T6472;
  wire[46:0] T6473;
  wire[46:0] T6474;
  wire[46:0] twiddle4_3_468_imag;
  wire[46:0] T6475;
  wire[46:0] T6476;
  wire[46:0] T6477;
  wire[45:0] T6478;
  wire[45:0] T6479;
  wire T6480;
  wire[46:0] twiddle4_3_469_imag;
  wire[46:0] T6481;
  wire[46:0] T6482;
  wire[46:0] T6483;
  wire[45:0] T6484;
  wire[45:0] T6485;
  wire T6486;
  wire T6487;
  wire[46:0] T6488;
  wire[46:0] twiddle4_3_470_imag;
  wire[46:0] T6489;
  wire[46:0] T6490;
  wire[46:0] T6491;
  wire[45:0] T6492;
  wire[45:0] T6493;
  wire T6494;
  wire[46:0] twiddle4_3_471_imag;
  wire[46:0] T6495;
  wire[46:0] T6496;
  wire[46:0] T6497;
  wire[45:0] T6498;
  wire[45:0] T6499;
  wire T6500;
  wire T6501;
  wire T6502;
  wire T6503;
  wire[46:0] T6504;
  wire[46:0] T6505;
  wire[46:0] T6506;
  wire[46:0] twiddle4_3_472_imag;
  wire[46:0] T6507;
  wire[46:0] T6508;
  wire[46:0] T6509;
  wire[45:0] T6510;
  wire[45:0] T6511;
  wire T6512;
  wire[46:0] twiddle4_3_473_imag;
  wire[46:0] T6513;
  wire[46:0] T6514;
  wire[46:0] T6515;
  wire[45:0] T6516;
  wire[45:0] T6517;
  wire T6518;
  wire T6519;
  wire[46:0] T6520;
  wire[46:0] twiddle4_3_474_imag;
  wire[46:0] T6521;
  wire[46:0] T6522;
  wire[46:0] T6523;
  wire[45:0] T6524;
  wire[45:0] T6525;
  wire T6526;
  wire[46:0] twiddle4_3_475_imag;
  wire[46:0] T6527;
  wire[46:0] T6528;
  wire[46:0] T6529;
  wire[45:0] T6530;
  wire[45:0] T6531;
  wire T6532;
  wire T6533;
  wire T6534;
  wire[46:0] T6535;
  wire[46:0] T6536;
  wire[46:0] twiddle4_3_476_imag;
  wire[46:0] T6537;
  wire[46:0] T6538;
  wire[46:0] T6539;
  wire[45:0] T6540;
  wire[45:0] T6541;
  wire T6542;
  wire[46:0] twiddle4_3_477_imag;
  wire[46:0] T6543;
  wire[46:0] T6544;
  wire[46:0] T6545;
  wire[45:0] T6546;
  wire[45:0] T6547;
  wire T6548;
  wire T6549;
  wire[46:0] T6550;
  wire[46:0] twiddle4_3_478_imag;
  wire[46:0] T6551;
  wire[46:0] T6552;
  wire[46:0] T6553;
  wire[45:0] T6554;
  wire[45:0] T6555;
  wire T6556;
  wire[46:0] twiddle4_3_479_imag;
  wire[46:0] T6557;
  wire[46:0] T6558;
  wire[46:0] T6559;
  wire[45:0] T6560;
  wire[45:0] T6561;
  wire T6562;
  wire T6563;
  wire T6564;
  wire T6565;
  wire T6566;
  wire T6567;
  wire[46:0] T6568;
  wire[46:0] T6569;
  wire[46:0] T6570;
  wire[46:0] T6571;
  wire[46:0] T6572;
  wire[46:0] twiddle4_3_480_imag;
  wire[46:0] T6573;
  wire[46:0] T6574;
  wire[46:0] T6575;
  wire[45:0] T6576;
  wire[45:0] T6577;
  wire T6578;
  wire[46:0] twiddle4_3_481_imag;
  wire[46:0] T6579;
  wire[46:0] T6580;
  wire[46:0] T6581;
  wire[45:0] T6582;
  wire[45:0] T6583;
  wire T6584;
  wire T6585;
  wire[46:0] T6586;
  wire[46:0] twiddle4_3_482_imag;
  wire[46:0] T6587;
  wire[46:0] T6588;
  wire[46:0] T6589;
  wire[45:0] T6590;
  wire[45:0] T6591;
  wire T6592;
  wire[46:0] twiddle4_3_483_imag;
  wire[46:0] T6593;
  wire[46:0] T6594;
  wire[46:0] T6595;
  wire[45:0] T6596;
  wire[45:0] T6597;
  wire T6598;
  wire T6599;
  wire T6600;
  wire[46:0] T6601;
  wire[46:0] T6602;
  wire[46:0] twiddle4_3_484_imag;
  wire[46:0] T6603;
  wire[46:0] T6604;
  wire[46:0] T6605;
  wire[45:0] T6606;
  wire[45:0] T6607;
  wire T6608;
  wire[46:0] twiddle4_3_485_imag;
  wire[46:0] T6609;
  wire[46:0] T6610;
  wire[46:0] T6611;
  wire[44:0] T6612;
  wire[44:0] T6613;
  wire[1:0] T6614;
  wire T6615;
  wire T6616;
  wire[46:0] T6617;
  wire[46:0] twiddle4_3_486_imag;
  wire[46:0] T6618;
  wire[46:0] T6619;
  wire[46:0] T6620;
  wire[44:0] T6621;
  wire[44:0] T6622;
  wire[1:0] T6623;
  wire T6624;
  wire[46:0] twiddle4_3_487_imag;
  wire[46:0] T6625;
  wire[46:0] T6626;
  wire[46:0] T6627;
  wire[44:0] T6628;
  wire[44:0] T6629;
  wire[1:0] T6630;
  wire T6631;
  wire T6632;
  wire T6633;
  wire T6634;
  wire[46:0] T6635;
  wire[46:0] T6636;
  wire[46:0] T6637;
  wire[46:0] twiddle4_3_488_imag;
  wire[46:0] T6638;
  wire[46:0] T6639;
  wire[46:0] T6640;
  wire[44:0] T6641;
  wire[44:0] T6642;
  wire[1:0] T6643;
  wire T6644;
  wire[46:0] twiddle4_3_489_imag;
  wire[46:0] T6645;
  wire[46:0] T6646;
  wire[46:0] T6647;
  wire[44:0] T6648;
  wire[44:0] T6649;
  wire[1:0] T6650;
  wire T6651;
  wire T6652;
  wire[46:0] T6653;
  wire[46:0] twiddle4_3_490_imag;
  wire[46:0] T6654;
  wire[46:0] T6655;
  wire[46:0] T6656;
  wire[44:0] T6657;
  wire[44:0] T6658;
  wire[1:0] T6659;
  wire T6660;
  wire[46:0] twiddle4_3_491_imag;
  wire[46:0] T6661;
  wire[46:0] T6662;
  wire[46:0] T6663;
  wire[44:0] T6664;
  wire[44:0] T6665;
  wire[1:0] T6666;
  wire T6667;
  wire T6668;
  wire T6669;
  wire[46:0] T6670;
  wire[46:0] T6671;
  wire[46:0] twiddle4_3_492_imag;
  wire[46:0] T6672;
  wire[46:0] T6673;
  wire[46:0] T6674;
  wire[44:0] T6675;
  wire[44:0] T6676;
  wire[1:0] T6677;
  wire T6678;
  wire[46:0] twiddle4_3_493_imag;
  wire[46:0] T6679;
  wire[46:0] T6680;
  wire[46:0] T6681;
  wire[44:0] T6682;
  wire[44:0] T6683;
  wire[1:0] T6684;
  wire T6685;
  wire T6686;
  wire[46:0] T6687;
  wire[46:0] twiddle4_3_494_imag;
  wire[46:0] T6688;
  wire[46:0] T6689;
  wire[46:0] T6690;
  wire[44:0] T6691;
  wire[44:0] T6692;
  wire[1:0] T6693;
  wire T6694;
  wire[46:0] twiddle4_3_495_imag;
  wire[46:0] T6695;
  wire[46:0] T6696;
  wire[46:0] T6697;
  wire[44:0] T6698;
  wire[44:0] T6699;
  wire[1:0] T6700;
  wire T6701;
  wire T6702;
  wire T6703;
  wire T6704;
  wire T6705;
  wire[46:0] T6706;
  wire[46:0] T6707;
  wire[46:0] T6708;
  wire[46:0] T6709;
  wire[46:0] twiddle4_3_496_imag;
  wire[46:0] T6710;
  wire[46:0] T6711;
  wire[46:0] T6712;
  wire[44:0] T6713;
  wire[44:0] T6714;
  wire[1:0] T6715;
  wire T6716;
  wire[46:0] twiddle4_3_497_imag;
  wire[46:0] T6717;
  wire[46:0] T6718;
  wire[46:0] T6719;
  wire[44:0] T6720;
  wire[44:0] T6721;
  wire[1:0] T6722;
  wire T6723;
  wire T6724;
  wire[46:0] T6725;
  wire[46:0] twiddle4_3_498_imag;
  wire[46:0] T6726;
  wire[46:0] T6727;
  wire[46:0] T6728;
  wire[44:0] T6729;
  wire[44:0] T6730;
  wire[1:0] T6731;
  wire T6732;
  wire[46:0] twiddle4_3_499_imag;
  wire[46:0] T6733;
  wire[46:0] T6734;
  wire[46:0] T6735;
  wire[43:0] T6736;
  wire[43:0] T6737;
  wire[2:0] T6738;
  wire T6739;
  wire T6740;
  wire T6741;
  wire[46:0] T6742;
  wire[46:0] T6743;
  wire[46:0] twiddle4_3_500_imag;
  wire[46:0] T6744;
  wire[46:0] T6745;
  wire[46:0] T6746;
  wire[43:0] T6747;
  wire[43:0] T6748;
  wire[2:0] T6749;
  wire T6750;
  wire[46:0] twiddle4_3_501_imag;
  wire[46:0] T6751;
  wire[46:0] T6752;
  wire[46:0] T6753;
  wire[43:0] T6754;
  wire[43:0] T6755;
  wire[2:0] T6756;
  wire T6757;
  wire T6758;
  wire[46:0] T6759;
  wire[46:0] twiddle4_3_502_imag;
  wire[46:0] T6760;
  wire[46:0] T6761;
  wire[46:0] T6762;
  wire[43:0] T6763;
  wire[43:0] T6764;
  wire[2:0] T6765;
  wire T6766;
  wire[46:0] twiddle4_3_503_imag;
  wire[46:0] T6767;
  wire[46:0] T6768;
  wire[46:0] T6769;
  wire[43:0] T6770;
  wire[43:0] T6771;
  wire[2:0] T6772;
  wire T6773;
  wire T6774;
  wire T6775;
  wire T6776;
  wire[46:0] T6777;
  wire[46:0] T6778;
  wire[46:0] T6779;
  wire[46:0] twiddle4_3_504_imag;
  wire[46:0] T6780;
  wire[46:0] T6781;
  wire[46:0] T6782;
  wire[43:0] T6783;
  wire[43:0] T6784;
  wire[2:0] T6785;
  wire T6786;
  wire[46:0] twiddle4_3_505_imag;
  wire[46:0] T6787;
  wire[46:0] T6788;
  wire[46:0] T6789;
  wire[43:0] T6790;
  wire[43:0] T6791;
  wire[2:0] T6792;
  wire T6793;
  wire T6794;
  wire[46:0] T6795;
  wire[46:0] twiddle4_3_506_imag;
  wire[46:0] T6796;
  wire[46:0] T6797;
  wire[46:0] T6798;
  wire[42:0] T6799;
  wire[42:0] T6800;
  wire[3:0] T6801;
  wire T6802;
  wire[46:0] twiddle4_3_507_imag;
  wire[46:0] T6803;
  wire[46:0] T6804;
  wire[46:0] T6805;
  wire[42:0] T6806;
  wire[42:0] T6807;
  wire[3:0] T6808;
  wire T6809;
  wire T6810;
  wire T6811;
  wire[46:0] T6812;
  wire[46:0] T6813;
  wire[46:0] twiddle4_3_508_imag;
  wire[46:0] T6814;
  wire[46:0] T6815;
  wire[46:0] T6816;
  wire[42:0] T6817;
  wire[42:0] T6818;
  wire[3:0] T6819;
  wire T6820;
  wire[46:0] twiddle4_3_509_imag;
  wire[46:0] T6821;
  wire[46:0] T6822;
  wire[46:0] T6823;
  wire[41:0] T6824;
  wire[41:0] T6825;
  wire[4:0] T6826;
  wire T6827;
  wire T6828;
  wire[46:0] T6829;
  wire[46:0] twiddle4_3_510_imag;
  wire[46:0] T6830;
  wire[46:0] T6831;
  wire[46:0] T6832;
  wire[41:0] T6833;
  wire[41:0] T6834;
  wire[4:0] T6835;
  wire T6836;
  wire[46:0] twiddle4_3_511_imag;
  wire[46:0] T6837;
  wire[46:0] T6838;
  wire[46:0] T6839;
  wire[40:0] T6840;
  wire[40:0] T6841;
  wire[5:0] T6842;
  wire T6843;
  wire T6844;
  wire T6845;
  wire T6846;
  wire T6847;
  wire T6848;
  wire T6849;
  wire T6850;
  wire T6851;
  wire T6852;
  wire T6853;
  wire[15:0] T6854;
  wire[47:0] T6855;
  wire[47:0] T6856;
  wire[47:0] T6857;
  wire[47:0] T6858;
  wire[47:0] T6859;
  wire[47:0] T6860;
  wire[47:0] T6861;
  wire[47:0] T6862;
  wire[47:0] T6863;
  wire[47:0] twiddle4_3_0_real;
  wire[47:0] T6864;
  wire[16:0] T6865;
  wire[16:0] T6866;
  wire[30:0] T6867;
  wire T6868;
  wire[47:0] T6869;
  wire[47:0] T6870;
  wire[47:0] T6871;
  wire[46:0] twiddle4_3_1_real;
  wire[46:0] T6872;
  wire[40:0] T6873;
  wire[40:0] T6874;
  wire[5:0] T6875;
  wire T6876;
  wire[46:0] T6877;
  wire[46:0] T6878;
  wire T6879;
  wire T6880;
  wire[47:0] T6881;
  wire[46:0] T6882;
  wire[46:0] twiddle4_3_2_real;
  wire[46:0] T6883;
  wire[41:0] T6884;
  wire[41:0] T6885;
  wire[4:0] T6886;
  wire T6887;
  wire[46:0] T6888;
  wire[46:0] T6889;
  wire[46:0] twiddle4_3_3_real;
  wire[46:0] T6890;
  wire[41:0] T6891;
  wire[41:0] T6892;
  wire[4:0] T6893;
  wire T6894;
  wire[46:0] T6895;
  wire[46:0] T6896;
  wire T6897;
  wire T6898;
  wire T6899;
  wire[47:0] T6900;
  wire[46:0] T6901;
  wire[46:0] T6902;
  wire[46:0] twiddle4_3_4_real;
  wire[46:0] T6903;
  wire[42:0] T6904;
  wire[42:0] T6905;
  wire[3:0] T6906;
  wire T6907;
  wire[46:0] T6908;
  wire[46:0] T6909;
  wire[46:0] twiddle4_3_5_real;
  wire[46:0] T6910;
  wire[42:0] T6911;
  wire[42:0] T6912;
  wire[3:0] T6913;
  wire T6914;
  wire[46:0] T6915;
  wire[46:0] T6916;
  wire T6917;
  wire[46:0] T6918;
  wire[46:0] twiddle4_3_6_real;
  wire[46:0] T6919;
  wire[42:0] T6920;
  wire[42:0] T6921;
  wire[3:0] T6922;
  wire T6923;
  wire[46:0] T6924;
  wire[46:0] T6925;
  wire[46:0] twiddle4_3_7_real;
  wire[46:0] T6926;
  wire[43:0] T6927;
  wire[43:0] T6928;
  wire[2:0] T6929;
  wire T6930;
  wire[46:0] T6931;
  wire[46:0] T6932;
  wire T6933;
  wire T6934;
  wire T6935;
  wire T6936;
  wire[47:0] T6937;
  wire[46:0] T6938;
  wire[46:0] T6939;
  wire[46:0] T6940;
  wire[46:0] twiddle4_3_8_real;
  wire[46:0] T6941;
  wire[43:0] T6942;
  wire[43:0] T6943;
  wire[2:0] T6944;
  wire T6945;
  wire[46:0] T6946;
  wire[46:0] T6947;
  wire[46:0] twiddle4_3_9_real;
  wire[46:0] T6948;
  wire[43:0] T6949;
  wire[43:0] T6950;
  wire[2:0] T6951;
  wire T6952;
  wire[46:0] T6953;
  wire[46:0] T6954;
  wire T6955;
  wire[46:0] T6956;
  wire[46:0] twiddle4_3_10_real;
  wire[46:0] T6957;
  wire[43:0] T6958;
  wire[43:0] T6959;
  wire[2:0] T6960;
  wire T6961;
  wire[46:0] T6962;
  wire[46:0] T6963;
  wire[46:0] twiddle4_3_11_real;
  wire[46:0] T6964;
  wire[43:0] T6965;
  wire[43:0] T6966;
  wire[2:0] T6967;
  wire T6968;
  wire[46:0] T6969;
  wire[46:0] T6970;
  wire T6971;
  wire T6972;
  wire[46:0] T6973;
  wire[46:0] T6974;
  wire[46:0] twiddle4_3_12_real;
  wire[46:0] T6975;
  wire[43:0] T6976;
  wire[43:0] T6977;
  wire[2:0] T6978;
  wire T6979;
  wire[46:0] T6980;
  wire[46:0] T6981;
  wire[46:0] twiddle4_3_13_real;
  wire[46:0] T6982;
  wire[43:0] T6983;
  wire[43:0] T6984;
  wire[2:0] T6985;
  wire T6986;
  wire[46:0] T6987;
  wire[46:0] T6988;
  wire T6989;
  wire[46:0] T6990;
  wire[46:0] twiddle4_3_14_real;
  wire[46:0] T6991;
  wire[44:0] T6992;
  wire[44:0] T6993;
  wire[1:0] T6994;
  wire T6995;
  wire[46:0] T6996;
  wire[46:0] T6997;
  wire[46:0] twiddle4_3_15_real;
  wire[46:0] T6998;
  wire[44:0] T6999;
  wire[44:0] T7000;
  wire[1:0] T7001;
  wire T7002;
  wire[46:0] T7003;
  wire[46:0] T7004;
  wire T7005;
  wire T7006;
  wire T7007;
  wire T7008;
  wire T7009;
  wire[47:0] T7010;
  wire[46:0] T7011;
  wire[46:0] T7012;
  wire[46:0] T7013;
  wire[46:0] T7014;
  wire[46:0] twiddle4_3_16_real;
  wire[46:0] T7015;
  wire[44:0] T7016;
  wire[44:0] T7017;
  wire[1:0] T7018;
  wire T7019;
  wire[46:0] T7020;
  wire[46:0] T7021;
  wire[46:0] twiddle4_3_17_real;
  wire[46:0] T7022;
  wire[44:0] T7023;
  wire[44:0] T7024;
  wire[1:0] T7025;
  wire T7026;
  wire[46:0] T7027;
  wire[46:0] T7028;
  wire T7029;
  wire[46:0] T7030;
  wire[46:0] twiddle4_3_18_real;
  wire[46:0] T7031;
  wire[44:0] T7032;
  wire[44:0] T7033;
  wire[1:0] T7034;
  wire T7035;
  wire[46:0] T7036;
  wire[46:0] T7037;
  wire[46:0] twiddle4_3_19_real;
  wire[46:0] T7038;
  wire[44:0] T7039;
  wire[44:0] T7040;
  wire[1:0] T7041;
  wire T7042;
  wire[46:0] T7043;
  wire[46:0] T7044;
  wire T7045;
  wire T7046;
  wire[46:0] T7047;
  wire[46:0] T7048;
  wire[46:0] twiddle4_3_20_real;
  wire[46:0] T7049;
  wire[44:0] T7050;
  wire[44:0] T7051;
  wire[1:0] T7052;
  wire T7053;
  wire[46:0] T7054;
  wire[46:0] T7055;
  wire[46:0] twiddle4_3_21_real;
  wire[46:0] T7056;
  wire[44:0] T7057;
  wire[44:0] T7058;
  wire[1:0] T7059;
  wire T7060;
  wire[46:0] T7061;
  wire[46:0] T7062;
  wire T7063;
  wire[46:0] T7064;
  wire[46:0] twiddle4_3_22_real;
  wire[46:0] T7065;
  wire[44:0] T7066;
  wire[44:0] T7067;
  wire[1:0] T7068;
  wire T7069;
  wire[46:0] T7070;
  wire[46:0] T7071;
  wire[46:0] twiddle4_3_23_real;
  wire[46:0] T7072;
  wire[44:0] T7073;
  wire[44:0] T7074;
  wire[1:0] T7075;
  wire T7076;
  wire[46:0] T7077;
  wire[46:0] T7078;
  wire T7079;
  wire T7080;
  wire T7081;
  wire[46:0] T7082;
  wire[46:0] T7083;
  wire[46:0] T7084;
  wire[46:0] twiddle4_3_24_real;
  wire[46:0] T7085;
  wire[44:0] T7086;
  wire[44:0] T7087;
  wire[1:0] T7088;
  wire T7089;
  wire[46:0] T7090;
  wire[46:0] T7091;
  wire[46:0] twiddle4_3_25_real;
  wire[46:0] T7092;
  wire[44:0] T7093;
  wire[44:0] T7094;
  wire[1:0] T7095;
  wire T7096;
  wire[46:0] T7097;
  wire[46:0] T7098;
  wire T7099;
  wire[46:0] T7100;
  wire[46:0] twiddle4_3_26_real;
  wire[46:0] T7101;
  wire[44:0] T7102;
  wire[44:0] T7103;
  wire[1:0] T7104;
  wire T7105;
  wire[46:0] T7106;
  wire[46:0] T7107;
  wire[46:0] twiddle4_3_27_real;
  wire[46:0] T7108;
  wire[44:0] T7109;
  wire[44:0] T7110;
  wire[1:0] T7111;
  wire T7112;
  wire[46:0] T7113;
  wire[46:0] T7114;
  wire T7115;
  wire T7116;
  wire[46:0] T7117;
  wire[46:0] T7118;
  wire[46:0] twiddle4_3_28_real;
  wire[46:0] T7119;
  wire[45:0] T7120;
  wire[45:0] T7121;
  wire T7122;
  wire[46:0] T7123;
  wire[46:0] T7124;
  wire[46:0] twiddle4_3_29_real;
  wire[46:0] T7125;
  wire[45:0] T7126;
  wire[45:0] T7127;
  wire T7128;
  wire[46:0] T7129;
  wire[46:0] T7130;
  wire T7131;
  wire[46:0] T7132;
  wire[46:0] twiddle4_3_30_real;
  wire[46:0] T7133;
  wire[45:0] T7134;
  wire[45:0] T7135;
  wire T7136;
  wire[46:0] T7137;
  wire[46:0] T7138;
  wire[46:0] twiddle4_3_31_real;
  wire[46:0] T7139;
  wire[45:0] T7140;
  wire[45:0] T7141;
  wire T7142;
  wire[46:0] T7143;
  wire[46:0] T7144;
  wire T7145;
  wire T7146;
  wire T7147;
  wire T7148;
  wire T7149;
  wire T7150;
  wire[47:0] T7151;
  wire[46:0] T7152;
  wire[46:0] T7153;
  wire[46:0] T7154;
  wire[46:0] T7155;
  wire[46:0] T7156;
  wire[46:0] twiddle4_3_32_real;
  wire[46:0] T7157;
  wire[45:0] T7158;
  wire[45:0] T7159;
  wire T7160;
  wire[46:0] T7161;
  wire[46:0] T7162;
  wire[46:0] twiddle4_3_33_real;
  wire[46:0] T7163;
  wire[45:0] T7164;
  wire[45:0] T7165;
  wire T7166;
  wire[46:0] T7167;
  wire[46:0] T7168;
  wire T7169;
  wire[46:0] T7170;
  wire[46:0] twiddle4_3_34_real;
  wire[46:0] T7171;
  wire[45:0] T7172;
  wire[45:0] T7173;
  wire T7174;
  wire[46:0] T7175;
  wire[46:0] T7176;
  wire[46:0] twiddle4_3_35_real;
  wire[46:0] T7177;
  wire[45:0] T7178;
  wire[45:0] T7179;
  wire T7180;
  wire[46:0] T7181;
  wire[46:0] T7182;
  wire T7183;
  wire T7184;
  wire[46:0] T7185;
  wire[46:0] T7186;
  wire[46:0] twiddle4_3_36_real;
  wire[46:0] T7187;
  wire[45:0] T7188;
  wire[45:0] T7189;
  wire T7190;
  wire[46:0] T7191;
  wire[46:0] T7192;
  wire[46:0] twiddle4_3_37_real;
  wire[46:0] T7193;
  wire[45:0] T7194;
  wire[45:0] T7195;
  wire T7196;
  wire[46:0] T7197;
  wire[46:0] T7198;
  wire T7199;
  wire[46:0] T7200;
  wire[46:0] twiddle4_3_38_real;
  wire[46:0] T7201;
  wire[45:0] T7202;
  wire[45:0] T7203;
  wire T7204;
  wire[46:0] T7205;
  wire[46:0] T7206;
  wire[46:0] twiddle4_3_39_real;
  wire[46:0] T7207;
  wire[45:0] T7208;
  wire[45:0] T7209;
  wire T7210;
  wire[46:0] T7211;
  wire[46:0] T7212;
  wire T7213;
  wire T7214;
  wire T7215;
  wire[46:0] T7216;
  wire[46:0] T7217;
  wire[46:0] T7218;
  wire[46:0] twiddle4_3_40_real;
  wire[46:0] T7219;
  wire[45:0] T7220;
  wire[45:0] T7221;
  wire T7222;
  wire[46:0] T7223;
  wire[46:0] T7224;
  wire[46:0] twiddle4_3_41_real;
  wire[46:0] T7225;
  wire[45:0] T7226;
  wire[45:0] T7227;
  wire T7228;
  wire[46:0] T7229;
  wire[46:0] T7230;
  wire T7231;
  wire[46:0] T7232;
  wire[46:0] twiddle4_3_42_real;
  wire[46:0] T7233;
  wire[45:0] T7234;
  wire[45:0] T7235;
  wire T7236;
  wire[46:0] T7237;
  wire[46:0] T7238;
  wire[46:0] twiddle4_3_43_real;
  wire[46:0] T7239;
  wire[45:0] T7240;
  wire[45:0] T7241;
  wire T7242;
  wire[46:0] T7243;
  wire[46:0] T7244;
  wire T7245;
  wire T7246;
  wire[46:0] T7247;
  wire[46:0] T7248;
  wire[46:0] twiddle4_3_44_real;
  wire[46:0] T7249;
  wire[45:0] T7250;
  wire[45:0] T7251;
  wire T7252;
  wire[46:0] T7253;
  wire[46:0] T7254;
  wire[46:0] twiddle4_3_45_real;
  wire[46:0] T7255;
  wire[45:0] T7256;
  wire[45:0] T7257;
  wire T7258;
  wire[46:0] T7259;
  wire[46:0] T7260;
  wire T7261;
  wire[46:0] T7262;
  wire[46:0] twiddle4_3_46_real;
  wire[46:0] T7263;
  wire[45:0] T7264;
  wire[45:0] T7265;
  wire T7266;
  wire[46:0] T7267;
  wire[46:0] T7268;
  wire[46:0] twiddle4_3_47_real;
  wire[46:0] T7269;
  wire[45:0] T7270;
  wire[45:0] T7271;
  wire T7272;
  wire[46:0] T7273;
  wire[46:0] T7274;
  wire T7275;
  wire T7276;
  wire T7277;
  wire T7278;
  wire[46:0] T7279;
  wire[46:0] T7280;
  wire[46:0] T7281;
  wire[46:0] T7282;
  wire[46:0] twiddle4_3_48_real;
  wire[46:0] T7283;
  wire[45:0] T7284;
  wire[45:0] T7285;
  wire T7286;
  wire[46:0] T7287;
  wire[46:0] T7288;
  wire[46:0] twiddle4_3_49_real;
  wire[46:0] T7289;
  wire[45:0] T7290;
  wire[45:0] T7291;
  wire T7292;
  wire[46:0] T7293;
  wire[46:0] T7294;
  wire T7295;
  wire[46:0] T7296;
  wire[46:0] twiddle4_3_50_real;
  wire[46:0] T7297;
  wire[45:0] T7298;
  wire[45:0] T7299;
  wire T7300;
  wire[46:0] T7301;
  wire[46:0] T7302;
  wire[46:0] twiddle4_3_51_real;
  wire[46:0] T7303;
  wire[45:0] T7304;
  wire[45:0] T7305;
  wire T7306;
  wire[46:0] T7307;
  wire[46:0] T7308;
  wire T7309;
  wire T7310;
  wire[46:0] T7311;
  wire[46:0] T7312;
  wire[46:0] twiddle4_3_52_real;
  wire[46:0] T7313;
  wire[45:0] T7314;
  wire[45:0] T7315;
  wire T7316;
  wire[46:0] T7317;
  wire[46:0] T7318;
  wire[46:0] twiddle4_3_53_real;
  wire[46:0] T7319;
  wire[45:0] T7320;
  wire[45:0] T7321;
  wire T7322;
  wire[46:0] T7323;
  wire[46:0] T7324;
  wire T7325;
  wire[46:0] T7326;
  wire[46:0] twiddle4_3_54_real;
  wire[46:0] T7327;
  wire[45:0] T7328;
  wire[45:0] T7329;
  wire T7330;
  wire[46:0] T7331;
  wire[46:0] T7332;
  wire[46:0] twiddle4_3_55_real;
  wire[46:0] T7333;
  wire[45:0] T7334;
  wire[45:0] T7335;
  wire T7336;
  wire[46:0] T7337;
  wire[46:0] T7338;
  wire T7339;
  wire T7340;
  wire T7341;
  wire[46:0] T7342;
  wire[46:0] T7343;
  wire[46:0] T7344;
  wire[46:0] twiddle4_3_56_real;
  wire[46:0] T7345;
  wire[45:0] T7346;
  wire[45:0] T7347;
  wire T7348;
  wire[46:0] T7349;
  wire[46:0] T7350;
  wire[46:0] twiddle4_3_57_real;
  wire[46:0] T7351;
  wire[46:0] T7352;
  wire[46:0] T7353;
  wire[46:0] T7354;
  wire T7355;
  wire[46:0] T7356;
  wire[46:0] twiddle4_3_58_real;
  wire[46:0] T7357;
  wire[46:0] T7358;
  wire[46:0] T7359;
  wire[46:0] T7360;
  wire[46:0] twiddle4_3_59_real;
  wire[46:0] T7361;
  wire[46:0] T7362;
  wire[46:0] T7363;
  wire[46:0] T7364;
  wire T7365;
  wire T7366;
  wire[46:0] T7367;
  wire[46:0] T7368;
  wire[46:0] twiddle4_3_60_real;
  wire[46:0] T7369;
  wire[46:0] T7370;
  wire[46:0] T7371;
  wire[46:0] T7372;
  wire[46:0] twiddle4_3_61_real;
  wire[46:0] T7373;
  wire[46:0] T7374;
  wire[46:0] T7375;
  wire[46:0] T7376;
  wire T7377;
  wire[46:0] T7378;
  wire[46:0] twiddle4_3_62_real;
  wire[46:0] T7379;
  wire[46:0] T7380;
  wire[46:0] T7381;
  wire[46:0] T7382;
  wire[46:0] twiddle4_3_63_real;
  wire[46:0] T7383;
  wire[46:0] T7384;
  wire[46:0] T7385;
  wire[46:0] T7386;
  wire T7387;
  wire T7388;
  wire T7389;
  wire T7390;
  wire T7391;
  wire T7392;
  wire T7393;
  wire[47:0] T7394;
  wire[46:0] T7395;
  wire[46:0] T7396;
  wire[46:0] T7397;
  wire[46:0] T7398;
  wire[46:0] T7399;
  wire[46:0] T7400;
  wire[46:0] twiddle4_3_64_real;
  wire[46:0] T7401;
  wire[46:0] T7402;
  wire[46:0] T7403;
  wire[46:0] T7404;
  wire[46:0] twiddle4_3_65_real;
  wire[46:0] T7405;
  wire[46:0] T7406;
  wire[46:0] T7407;
  wire[46:0] T7408;
  wire T7409;
  wire[46:0] T7410;
  wire[46:0] twiddle4_3_66_real;
  wire[46:0] T7411;
  wire[46:0] T7412;
  wire[46:0] T7413;
  wire[46:0] T7414;
  wire[46:0] twiddle4_3_67_real;
  wire[46:0] T7415;
  wire[46:0] T7416;
  wire[46:0] T7417;
  wire[46:0] T7418;
  wire T7419;
  wire T7420;
  wire[46:0] T7421;
  wire[46:0] T7422;
  wire[46:0] twiddle4_3_68_real;
  wire[46:0] T7423;
  wire[46:0] T7424;
  wire[46:0] T7425;
  wire[46:0] T7426;
  wire[46:0] twiddle4_3_69_real;
  wire[46:0] T7427;
  wire[46:0] T7428;
  wire[46:0] T7429;
  wire[46:0] T7430;
  wire T7431;
  wire[46:0] T7432;
  wire[46:0] twiddle4_3_70_real;
  wire[46:0] T7433;
  wire[46:0] T7434;
  wire[46:0] T7435;
  wire[46:0] T7436;
  wire[46:0] twiddle4_3_71_real;
  wire[46:0] T7437;
  wire[46:0] T7438;
  wire[46:0] T7439;
  wire[46:0] T7440;
  wire T7441;
  wire T7442;
  wire T7443;
  wire[46:0] T7444;
  wire[46:0] T7445;
  wire[46:0] T7446;
  wire[46:0] twiddle4_3_72_real;
  wire[46:0] T7447;
  wire[46:0] T7448;
  wire[46:0] T7449;
  wire[46:0] T7450;
  wire[46:0] twiddle4_3_73_real;
  wire[46:0] T7451;
  wire[46:0] T7452;
  wire[46:0] T7453;
  wire[46:0] T7454;
  wire T7455;
  wire[46:0] T7456;
  wire[46:0] twiddle4_3_74_real;
  wire[46:0] T7457;
  wire[46:0] T7458;
  wire[46:0] T7459;
  wire[46:0] T7460;
  wire[46:0] twiddle4_3_75_real;
  wire[46:0] T7461;
  wire[46:0] T7462;
  wire[46:0] T7463;
  wire[46:0] T7464;
  wire T7465;
  wire T7466;
  wire[46:0] T7467;
  wire[46:0] T7468;
  wire[46:0] twiddle4_3_76_real;
  wire[46:0] T7469;
  wire[46:0] T7470;
  wire[46:0] T7471;
  wire[46:0] T7472;
  wire[46:0] twiddle4_3_77_real;
  wire[46:0] T7473;
  wire[46:0] T7474;
  wire[46:0] T7475;
  wire[46:0] T7476;
  wire T7477;
  wire[46:0] T7478;
  wire[46:0] twiddle4_3_78_real;
  wire[46:0] T7479;
  wire[46:0] T7480;
  wire[46:0] T7481;
  wire[46:0] T7482;
  wire[46:0] twiddle4_3_79_real;
  wire[46:0] T7483;
  wire[46:0] T7484;
  wire[46:0] T7485;
  wire[46:0] T7486;
  wire T7487;
  wire T7488;
  wire T7489;
  wire T7490;
  wire[46:0] T7491;
  wire[46:0] T7492;
  wire[46:0] T7493;
  wire[46:0] T7494;
  wire[46:0] twiddle4_3_80_real;
  wire[46:0] T7495;
  wire[46:0] T7496;
  wire[46:0] T7497;
  wire[46:0] T7498;
  wire[46:0] twiddle4_3_81_real;
  wire[46:0] T7499;
  wire[46:0] T7500;
  wire[46:0] T7501;
  wire[46:0] T7502;
  wire T7503;
  wire[46:0] T7504;
  wire[46:0] twiddle4_3_82_real;
  wire[46:0] T7505;
  wire[46:0] T7506;
  wire[46:0] T7507;
  wire[46:0] T7508;
  wire[46:0] twiddle4_3_83_real;
  wire[46:0] T7509;
  wire[46:0] T7510;
  wire[46:0] T7511;
  wire[46:0] T7512;
  wire T7513;
  wire T7514;
  wire[46:0] T7515;
  wire[46:0] T7516;
  wire[46:0] twiddle4_3_84_real;
  wire[46:0] T7517;
  wire[46:0] T7518;
  wire[46:0] T7519;
  wire[46:0] T7520;
  wire[46:0] twiddle4_3_85_real;
  wire[46:0] T7521;
  wire[46:0] T7522;
  wire[46:0] T7523;
  wire[46:0] T7524;
  wire T7525;
  wire[46:0] T7526;
  wire[46:0] twiddle4_3_86_real;
  wire[46:0] T7527;
  wire[46:0] T7528;
  wire[46:0] T7529;
  wire[46:0] T7530;
  wire[46:0] twiddle4_3_87_real;
  wire[46:0] T7531;
  wire[46:0] T7532;
  wire[46:0] T7533;
  wire[46:0] T7534;
  wire T7535;
  wire T7536;
  wire T7537;
  wire[46:0] T7538;
  wire[46:0] T7539;
  wire[46:0] T7540;
  wire[46:0] twiddle4_3_88_real;
  wire[46:0] T7541;
  wire[46:0] T7542;
  wire[46:0] T7543;
  wire[46:0] T7544;
  wire[46:0] twiddle4_3_89_real;
  wire[46:0] T7545;
  wire[46:0] T7546;
  wire[46:0] T7547;
  wire[46:0] T7548;
  wire T7549;
  wire[46:0] T7550;
  wire[46:0] twiddle4_3_90_real;
  wire[46:0] T7551;
  wire[46:0] T7552;
  wire[46:0] T7553;
  wire[46:0] T7554;
  wire[46:0] twiddle4_3_91_real;
  wire[46:0] T7555;
  wire[46:0] T7556;
  wire[46:0] T7557;
  wire[46:0] T7558;
  wire T7559;
  wire T7560;
  wire[46:0] T7561;
  wire[46:0] T7562;
  wire[46:0] twiddle4_3_92_real;
  wire[46:0] T7563;
  wire[46:0] T7564;
  wire[46:0] T7565;
  wire[46:0] T7566;
  wire[46:0] twiddle4_3_93_real;
  wire[46:0] T7567;
  wire[46:0] T7568;
  wire[46:0] T7569;
  wire[46:0] T7570;
  wire T7571;
  wire[46:0] T7572;
  wire[46:0] twiddle4_3_94_real;
  wire[46:0] T7573;
  wire[46:0] T7574;
  wire[46:0] T7575;
  wire[46:0] T7576;
  wire[46:0] twiddle4_3_95_real;
  wire[46:0] T7577;
  wire[46:0] T7578;
  wire[46:0] T7579;
  wire[46:0] T7580;
  wire T7581;
  wire T7582;
  wire T7583;
  wire T7584;
  wire T7585;
  wire[46:0] T7586;
  wire[46:0] T7587;
  wire[46:0] T7588;
  wire[46:0] T7589;
  wire[46:0] T7590;
  wire[46:0] twiddle4_3_96_real;
  wire[46:0] T7591;
  wire[46:0] T7592;
  wire[46:0] T7593;
  wire[46:0] T7594;
  wire[46:0] twiddle4_3_97_real;
  wire[46:0] T7595;
  wire[46:0] T7596;
  wire[46:0] T7597;
  wire[46:0] T7598;
  wire T7599;
  wire[46:0] T7600;
  wire[46:0] twiddle4_3_98_real;
  wire[46:0] T7601;
  wire[46:0] T7602;
  wire[46:0] T7603;
  wire[46:0] T7604;
  wire[46:0] twiddle4_3_99_real;
  wire[46:0] T7605;
  wire[46:0] T7606;
  wire[46:0] T7607;
  wire[46:0] T7608;
  wire T7609;
  wire T7610;
  wire[46:0] T7611;
  wire[46:0] T7612;
  wire[46:0] twiddle4_3_100_real;
  wire[46:0] T7613;
  wire[46:0] T7614;
  wire[46:0] T7615;
  wire[46:0] T7616;
  wire[46:0] twiddle4_3_101_real;
  wire[46:0] T7617;
  wire[46:0] T7618;
  wire[46:0] T7619;
  wire[46:0] T7620;
  wire T7621;
  wire[46:0] T7622;
  wire[46:0] twiddle4_3_102_real;
  wire[46:0] T7623;
  wire[46:0] T7624;
  wire[46:0] T7625;
  wire[46:0] T7626;
  wire[46:0] twiddle4_3_103_real;
  wire[46:0] T7627;
  wire[46:0] T7628;
  wire[46:0] T7629;
  wire[46:0] T7630;
  wire T7631;
  wire T7632;
  wire T7633;
  wire[46:0] T7634;
  wire[46:0] T7635;
  wire[46:0] T7636;
  wire[46:0] twiddle4_3_104_real;
  wire[46:0] T7637;
  wire[46:0] T7638;
  wire[46:0] T7639;
  wire[46:0] T7640;
  wire[46:0] twiddle4_3_105_real;
  wire[46:0] T7641;
  wire[46:0] T7642;
  wire[46:0] T7643;
  wire[46:0] T7644;
  wire T7645;
  wire[46:0] T7646;
  wire[46:0] twiddle4_3_106_real;
  wire[46:0] T7647;
  wire[46:0] T7648;
  wire[46:0] T7649;
  wire[46:0] T7650;
  wire[46:0] twiddle4_3_107_real;
  wire[46:0] T7651;
  wire[46:0] T7652;
  wire[46:0] T7653;
  wire[46:0] T7654;
  wire T7655;
  wire T7656;
  wire[46:0] T7657;
  wire[46:0] T7658;
  wire[46:0] twiddle4_3_108_real;
  wire[46:0] T7659;
  wire[46:0] T7660;
  wire[46:0] T7661;
  wire[46:0] T7662;
  wire[46:0] twiddle4_3_109_real;
  wire[46:0] T7663;
  wire[46:0] T7664;
  wire[46:0] T7665;
  wire[46:0] T7666;
  wire T7667;
  wire[46:0] T7668;
  wire[46:0] twiddle4_3_110_real;
  wire[46:0] T7669;
  wire[46:0] T7670;
  wire[46:0] T7671;
  wire[46:0] T7672;
  wire[46:0] twiddle4_3_111_real;
  wire[46:0] T7673;
  wire[46:0] T7674;
  wire[46:0] T7675;
  wire[46:0] T7676;
  wire T7677;
  wire T7678;
  wire T7679;
  wire T7680;
  wire[46:0] T7681;
  wire[46:0] T7682;
  wire[46:0] T7683;
  wire[46:0] T7684;
  wire[46:0] twiddle4_3_112_real;
  wire[46:0] T7685;
  wire[46:0] T7686;
  wire[46:0] T7687;
  wire[46:0] T7688;
  wire[46:0] twiddle4_3_113_real;
  wire[46:0] T7689;
  wire[46:0] T7690;
  wire[46:0] T7691;
  wire[46:0] T7692;
  wire T7693;
  wire[46:0] T7694;
  wire[46:0] twiddle4_3_114_real;
  wire[46:0] T7695;
  wire[46:0] T7696;
  wire[46:0] T7697;
  wire[45:0] T7698;
  wire[45:0] T7699;
  wire T7700;
  wire[46:0] twiddle4_3_115_real;
  wire[46:0] T7701;
  wire[46:0] T7702;
  wire[46:0] T7703;
  wire[45:0] T7704;
  wire[45:0] T7705;
  wire T7706;
  wire T7707;
  wire T7708;
  wire[46:0] T7709;
  wire[46:0] T7710;
  wire[46:0] twiddle4_3_116_real;
  wire[46:0] T7711;
  wire[46:0] T7712;
  wire[46:0] T7713;
  wire[45:0] T7714;
  wire[45:0] T7715;
  wire T7716;
  wire[46:0] twiddle4_3_117_real;
  wire[46:0] T7717;
  wire[46:0] T7718;
  wire[46:0] T7719;
  wire[45:0] T7720;
  wire[45:0] T7721;
  wire T7722;
  wire T7723;
  wire[46:0] T7724;
  wire[46:0] twiddle4_3_118_real;
  wire[46:0] T7725;
  wire[46:0] T7726;
  wire[46:0] T7727;
  wire[45:0] T7728;
  wire[45:0] T7729;
  wire T7730;
  wire[46:0] twiddle4_3_119_real;
  wire[46:0] T7731;
  wire[46:0] T7732;
  wire[46:0] T7733;
  wire[45:0] T7734;
  wire[45:0] T7735;
  wire T7736;
  wire T7737;
  wire T7738;
  wire T7739;
  wire[46:0] T7740;
  wire[46:0] T7741;
  wire[46:0] T7742;
  wire[46:0] twiddle4_3_120_real;
  wire[46:0] T7743;
  wire[46:0] T7744;
  wire[46:0] T7745;
  wire[45:0] T7746;
  wire[45:0] T7747;
  wire T7748;
  wire[46:0] twiddle4_3_121_real;
  wire[46:0] T7749;
  wire[46:0] T7750;
  wire[46:0] T7751;
  wire[45:0] T7752;
  wire[45:0] T7753;
  wire T7754;
  wire T7755;
  wire[46:0] T7756;
  wire[46:0] twiddle4_3_122_real;
  wire[46:0] T7757;
  wire[46:0] T7758;
  wire[46:0] T7759;
  wire[45:0] T7760;
  wire[45:0] T7761;
  wire T7762;
  wire[46:0] twiddle4_3_123_real;
  wire[46:0] T7763;
  wire[46:0] T7764;
  wire[46:0] T7765;
  wire[45:0] T7766;
  wire[45:0] T7767;
  wire T7768;
  wire T7769;
  wire T7770;
  wire[46:0] T7771;
  wire[46:0] T7772;
  wire[46:0] twiddle4_3_124_real;
  wire[46:0] T7773;
  wire[46:0] T7774;
  wire[46:0] T7775;
  wire[45:0] T7776;
  wire[45:0] T7777;
  wire T7778;
  wire[46:0] twiddle4_3_125_real;
  wire[46:0] T7779;
  wire[46:0] T7780;
  wire[46:0] T7781;
  wire[45:0] T7782;
  wire[45:0] T7783;
  wire T7784;
  wire T7785;
  wire[46:0] T7786;
  wire[46:0] twiddle4_3_126_real;
  wire[46:0] T7787;
  wire[46:0] T7788;
  wire[46:0] T7789;
  wire[45:0] T7790;
  wire[45:0] T7791;
  wire T7792;
  wire[46:0] twiddle4_3_127_real;
  wire[46:0] T7793;
  wire[46:0] T7794;
  wire[46:0] T7795;
  wire[45:0] T7796;
  wire[45:0] T7797;
  wire T7798;
  wire T7799;
  wire T7800;
  wire T7801;
  wire T7802;
  wire T7803;
  wire T7804;
  wire T7805;
  wire T7806;
  wire[47:0] T7807;
  wire[46:0] T7808;
  wire[46:0] T7809;
  wire[46:0] T7810;
  wire[46:0] T7811;
  wire[46:0] T7812;
  wire[46:0] T7813;
  wire[46:0] T7814;
  wire[46:0] twiddle4_3_128_real;
  wire[46:0] T7815;
  wire[46:0] T7816;
  wire[46:0] T7817;
  wire[45:0] T7818;
  wire[45:0] T7819;
  wire T7820;
  wire[46:0] twiddle4_3_129_real;
  wire[46:0] T7821;
  wire[46:0] T7822;
  wire[46:0] T7823;
  wire[45:0] T7824;
  wire[45:0] T7825;
  wire T7826;
  wire T7827;
  wire[46:0] T7828;
  wire[46:0] twiddle4_3_130_real;
  wire[46:0] T7829;
  wire[46:0] T7830;
  wire[46:0] T7831;
  wire[45:0] T7832;
  wire[45:0] T7833;
  wire T7834;
  wire[46:0] twiddle4_3_131_real;
  wire[46:0] T7835;
  wire[46:0] T7836;
  wire[46:0] T7837;
  wire[45:0] T7838;
  wire[45:0] T7839;
  wire T7840;
  wire T7841;
  wire T7842;
  wire[46:0] T7843;
  wire[46:0] T7844;
  wire[46:0] twiddle4_3_132_real;
  wire[46:0] T7845;
  wire[46:0] T7846;
  wire[46:0] T7847;
  wire[45:0] T7848;
  wire[45:0] T7849;
  wire T7850;
  wire[46:0] twiddle4_3_133_real;
  wire[46:0] T7851;
  wire[46:0] T7852;
  wire[46:0] T7853;
  wire[45:0] T7854;
  wire[45:0] T7855;
  wire T7856;
  wire T7857;
  wire[46:0] T7858;
  wire[46:0] twiddle4_3_134_real;
  wire[46:0] T7859;
  wire[46:0] T7860;
  wire[46:0] T7861;
  wire[45:0] T7862;
  wire[45:0] T7863;
  wire T7864;
  wire[46:0] twiddle4_3_135_real;
  wire[46:0] T7865;
  wire[46:0] T7866;
  wire[46:0] T7867;
  wire[45:0] T7868;
  wire[45:0] T7869;
  wire T7870;
  wire T7871;
  wire T7872;
  wire T7873;
  wire[46:0] T7874;
  wire[46:0] T7875;
  wire[46:0] T7876;
  wire[46:0] twiddle4_3_136_real;
  wire[46:0] T7877;
  wire[46:0] T7878;
  wire[46:0] T7879;
  wire[45:0] T7880;
  wire[45:0] T7881;
  wire T7882;
  wire[46:0] twiddle4_3_137_real;
  wire[46:0] T7883;
  wire[46:0] T7884;
  wire[46:0] T7885;
  wire[45:0] T7886;
  wire[45:0] T7887;
  wire T7888;
  wire T7889;
  wire[46:0] T7890;
  wire[46:0] twiddle4_3_138_real;
  wire[46:0] T7891;
  wire[46:0] T7892;
  wire[46:0] T7893;
  wire[45:0] T7894;
  wire[45:0] T7895;
  wire T7896;
  wire[46:0] twiddle4_3_139_real;
  wire[46:0] T7897;
  wire[46:0] T7898;
  wire[46:0] T7899;
  wire[45:0] T7900;
  wire[45:0] T7901;
  wire T7902;
  wire T7903;
  wire T7904;
  wire[46:0] T7905;
  wire[46:0] T7906;
  wire[46:0] twiddle4_3_140_real;
  wire[46:0] T7907;
  wire[46:0] T7908;
  wire[46:0] T7909;
  wire[45:0] T7910;
  wire[45:0] T7911;
  wire T7912;
  wire[46:0] twiddle4_3_141_real;
  wire[46:0] T7913;
  wire[46:0] T7914;
  wire[46:0] T7915;
  wire[45:0] T7916;
  wire[45:0] T7917;
  wire T7918;
  wire T7919;
  wire[46:0] T7920;
  wire[46:0] twiddle4_3_142_real;
  wire[46:0] T7921;
  wire[46:0] T7922;
  wire[46:0] T7923;
  wire[45:0] T7924;
  wire[45:0] T7925;
  wire T7926;
  wire[46:0] twiddle4_3_143_real;
  wire[46:0] T7927;
  wire[46:0] T7928;
  wire[46:0] T7929;
  wire[45:0] T7930;
  wire[45:0] T7931;
  wire T7932;
  wire T7933;
  wire T7934;
  wire T7935;
  wire T7936;
  wire[46:0] T7937;
  wire[46:0] T7938;
  wire[46:0] T7939;
  wire[46:0] T7940;
  wire[46:0] twiddle4_3_144_real;
  wire[46:0] T7941;
  wire[46:0] T7942;
  wire[46:0] T7943;
  wire[44:0] T7944;
  wire[44:0] T7945;
  wire[1:0] T7946;
  wire T7947;
  wire[46:0] twiddle4_3_145_real;
  wire[46:0] T7948;
  wire[46:0] T7949;
  wire[46:0] T7950;
  wire[44:0] T7951;
  wire[44:0] T7952;
  wire[1:0] T7953;
  wire T7954;
  wire T7955;
  wire[46:0] T7956;
  wire[46:0] twiddle4_3_146_real;
  wire[46:0] T7957;
  wire[46:0] T7958;
  wire[46:0] T7959;
  wire[44:0] T7960;
  wire[44:0] T7961;
  wire[1:0] T7962;
  wire T7963;
  wire[46:0] twiddle4_3_147_real;
  wire[46:0] T7964;
  wire[46:0] T7965;
  wire[46:0] T7966;
  wire[44:0] T7967;
  wire[44:0] T7968;
  wire[1:0] T7969;
  wire T7970;
  wire T7971;
  wire T7972;
  wire[46:0] T7973;
  wire[46:0] T7974;
  wire[46:0] twiddle4_3_148_real;
  wire[46:0] T7975;
  wire[46:0] T7976;
  wire[46:0] T7977;
  wire[44:0] T7978;
  wire[44:0] T7979;
  wire[1:0] T7980;
  wire T7981;
  wire[46:0] twiddle4_3_149_real;
  wire[46:0] T7982;
  wire[46:0] T7983;
  wire[46:0] T7984;
  wire[44:0] T7985;
  wire[44:0] T7986;
  wire[1:0] T7987;
  wire T7988;
  wire T7989;
  wire[46:0] T7990;
  wire[46:0] twiddle4_3_150_real;
  wire[46:0] T7991;
  wire[46:0] T7992;
  wire[46:0] T7993;
  wire[44:0] T7994;
  wire[44:0] T7995;
  wire[1:0] T7996;
  wire T7997;
  wire[46:0] twiddle4_3_151_real;
  wire[46:0] T7998;
  wire[46:0] T7999;
  wire[46:0] T8000;
  wire[44:0] T8001;
  wire[44:0] T8002;
  wire[1:0] T8003;
  wire T8004;
  wire T8005;
  wire T8006;
  wire T8007;
  wire[46:0] T8008;
  wire[46:0] T8009;
  wire[46:0] T8010;
  wire[46:0] twiddle4_3_152_real;
  wire[46:0] T8011;
  wire[46:0] T8012;
  wire[46:0] T8013;
  wire[44:0] T8014;
  wire[44:0] T8015;
  wire[1:0] T8016;
  wire T8017;
  wire[46:0] twiddle4_3_153_real;
  wire[46:0] T8018;
  wire[46:0] T8019;
  wire[46:0] T8020;
  wire[44:0] T8021;
  wire[44:0] T8022;
  wire[1:0] T8023;
  wire T8024;
  wire T8025;
  wire[46:0] T8026;
  wire[46:0] twiddle4_3_154_real;
  wire[46:0] T8027;
  wire[46:0] T8028;
  wire[46:0] T8029;
  wire[44:0] T8030;
  wire[44:0] T8031;
  wire[1:0] T8032;
  wire T8033;
  wire[46:0] twiddle4_3_155_real;
  wire[46:0] T8034;
  wire[46:0] T8035;
  wire[46:0] T8036;
  wire[44:0] T8037;
  wire[44:0] T8038;
  wire[1:0] T8039;
  wire T8040;
  wire T8041;
  wire T8042;
  wire[46:0] T8043;
  wire[46:0] T8044;
  wire[46:0] twiddle4_3_156_real;
  wire[46:0] T8045;
  wire[46:0] T8046;
  wire[46:0] T8047;
  wire[44:0] T8048;
  wire[44:0] T8049;
  wire[1:0] T8050;
  wire T8051;
  wire[46:0] twiddle4_3_157_real;
  wire[46:0] T8052;
  wire[46:0] T8053;
  wire[46:0] T8054;
  wire[44:0] T8055;
  wire[44:0] T8056;
  wire[1:0] T8057;
  wire T8058;
  wire T8059;
  wire[46:0] T8060;
  wire[46:0] twiddle4_3_158_real;
  wire[46:0] T8061;
  wire[46:0] T8062;
  wire[46:0] T8063;
  wire[43:0] T8064;
  wire[43:0] T8065;
  wire[2:0] T8066;
  wire T8067;
  wire[46:0] twiddle4_3_159_real;
  wire[46:0] T8068;
  wire[46:0] T8069;
  wire[46:0] T8070;
  wire[43:0] T8071;
  wire[43:0] T8072;
  wire[2:0] T8073;
  wire T8074;
  wire T8075;
  wire T8076;
  wire T8077;
  wire T8078;
  wire T8079;
  wire[46:0] T8080;
  wire[46:0] T8081;
  wire[46:0] T8082;
  wire[46:0] T8083;
  wire[46:0] T8084;
  wire[46:0] twiddle4_3_160_real;
  wire[46:0] T8085;
  wire[46:0] T8086;
  wire[46:0] T8087;
  wire[43:0] T8088;
  wire[43:0] T8089;
  wire[2:0] T8090;
  wire T8091;
  wire[46:0] twiddle4_3_161_real;
  wire[46:0] T8092;
  wire[46:0] T8093;
  wire[46:0] T8094;
  wire[43:0] T8095;
  wire[43:0] T8096;
  wire[2:0] T8097;
  wire T8098;
  wire T8099;
  wire[46:0] T8100;
  wire[46:0] twiddle4_3_162_real;
  wire[46:0] T8101;
  wire[46:0] T8102;
  wire[46:0] T8103;
  wire[43:0] T8104;
  wire[43:0] T8105;
  wire[2:0] T8106;
  wire T8107;
  wire[46:0] twiddle4_3_163_real;
  wire[46:0] T8108;
  wire[46:0] T8109;
  wire[46:0] T8110;
  wire[43:0] T8111;
  wire[43:0] T8112;
  wire[2:0] T8113;
  wire T8114;
  wire T8115;
  wire T8116;
  wire[46:0] T8117;
  wire[46:0] T8118;
  wire[46:0] twiddle4_3_164_real;
  wire[46:0] T8119;
  wire[46:0] T8120;
  wire[46:0] T8121;
  wire[42:0] T8122;
  wire[42:0] T8123;
  wire[3:0] T8124;
  wire T8125;
  wire[46:0] twiddle4_3_165_real;
  wire[46:0] T8126;
  wire[46:0] T8127;
  wire[46:0] T8128;
  wire[42:0] T8129;
  wire[42:0] T8130;
  wire[3:0] T8131;
  wire T8132;
  wire T8133;
  wire[46:0] T8134;
  wire[46:0] twiddle4_3_166_real;
  wire[46:0] T8135;
  wire[46:0] T8136;
  wire[46:0] T8137;
  wire[42:0] T8138;
  wire[42:0] T8139;
  wire[3:0] T8140;
  wire T8141;
  wire[46:0] twiddle4_3_167_real;
  wire[46:0] T8142;
  wire[46:0] T8143;
  wire[46:0] T8144;
  wire[42:0] T8145;
  wire[42:0] T8146;
  wire[3:0] T8147;
  wire T8148;
  wire T8149;
  wire T8150;
  wire T8151;
  wire[46:0] T8152;
  wire[46:0] T8153;
  wire[46:0] T8154;
  wire[46:0] twiddle4_3_168_real;
  wire[46:0] T8155;
  wire[46:0] T8156;
  wire[46:0] T8157;
  wire[41:0] T8158;
  wire[41:0] T8159;
  wire[4:0] T8160;
  wire T8161;
  wire[46:0] twiddle4_3_169_real;
  wire[46:0] T8162;
  wire[46:0] T8163;
  wire[46:0] T8164;
  wire[40:0] T8165;
  wire[40:0] T8166;
  wire[5:0] T8167;
  wire T8168;
  wire T8169;
  wire[46:0] T8170;
  wire[46:0] twiddle4_3_170_real;
  wire[46:0] T8171;
  wire[46:0] T8172;
  wire[46:0] T8173;
  wire[39:0] T8174;
  wire[39:0] T8175;
  wire[6:0] T8176;
  wire T8177;
  wire[46:0] twiddle4_3_171_real;
  wire[46:0] T8178;
  wire[46:0] T8179;
  wire[46:0] T8180;
  wire[38:0] T8181;
  wire[38:0] T8182;
  wire[7:0] T8183;
  wire T8184;
  wire T8185;
  wire T8186;
  wire[46:0] T8187;
  wire[46:0] T8188;
  wire[46:0] twiddle4_3_172_real;
  wire[46:0] T8189;
  wire[46:0] T8190;
  wire[46:0] T8191;
  wire[40:0] T8192;
  wire[40:0] T8193;
  wire[5:0] T8194;
  wire T8195;
  wire[46:0] twiddle4_3_173_real;
  wire[46:0] T8196;
  wire[46:0] T8197;
  wire[46:0] T8198;
  wire[41:0] T8199;
  wire[41:0] T8200;
  wire[4:0] T8201;
  wire T8202;
  wire T8203;
  wire[46:0] T8204;
  wire[46:0] twiddle4_3_174_real;
  wire[46:0] T8205;
  wire[46:0] T8206;
  wire[46:0] T8207;
  wire[41:0] T8208;
  wire[41:0] T8209;
  wire[4:0] T8210;
  wire T8211;
  wire[46:0] twiddle4_3_175_real;
  wire[46:0] T8212;
  wire[46:0] T8213;
  wire[46:0] T8214;
  wire[42:0] T8215;
  wire[42:0] T8216;
  wire[3:0] T8217;
  wire T8218;
  wire T8219;
  wire T8220;
  wire T8221;
  wire T8222;
  wire[46:0] T8223;
  wire[46:0] T8224;
  wire[46:0] T8225;
  wire[46:0] T8226;
  wire[46:0] twiddle4_3_176_real;
  wire[46:0] T8227;
  wire[46:0] T8228;
  wire[46:0] T8229;
  wire[42:0] T8230;
  wire[42:0] T8231;
  wire[3:0] T8232;
  wire T8233;
  wire[46:0] twiddle4_3_177_real;
  wire[46:0] T8234;
  wire[46:0] T8235;
  wire[46:0] T8236;
  wire[42:0] T8237;
  wire[42:0] T8238;
  wire[3:0] T8239;
  wire T8240;
  wire T8241;
  wire[46:0] T8242;
  wire[46:0] twiddle4_3_178_real;
  wire[46:0] T8243;
  wire[46:0] T8244;
  wire[46:0] T8245;
  wire[43:0] T8246;
  wire[43:0] T8247;
  wire[2:0] T8248;
  wire T8249;
  wire[46:0] twiddle4_3_179_real;
  wire[46:0] T8250;
  wire[46:0] T8251;
  wire[46:0] T8252;
  wire[43:0] T8253;
  wire[43:0] T8254;
  wire[2:0] T8255;
  wire T8256;
  wire T8257;
  wire T8258;
  wire[46:0] T8259;
  wire[46:0] T8260;
  wire[46:0] twiddle4_3_180_real;
  wire[46:0] T8261;
  wire[46:0] T8262;
  wire[46:0] T8263;
  wire[43:0] T8264;
  wire[43:0] T8265;
  wire[2:0] T8266;
  wire T8267;
  wire[46:0] twiddle4_3_181_real;
  wire[46:0] T8268;
  wire[46:0] T8269;
  wire[46:0] T8270;
  wire[43:0] T8271;
  wire[43:0] T8272;
  wire[2:0] T8273;
  wire T8274;
  wire T8275;
  wire[46:0] T8276;
  wire[46:0] twiddle4_3_182_real;
  wire[46:0] T8277;
  wire[46:0] T8278;
  wire[46:0] T8279;
  wire[43:0] T8280;
  wire[43:0] T8281;
  wire[2:0] T8282;
  wire T8283;
  wire[46:0] twiddle4_3_183_real;
  wire[46:0] T8284;
  wire[46:0] T8285;
  wire[46:0] T8286;
  wire[43:0] T8287;
  wire[43:0] T8288;
  wire[2:0] T8289;
  wire T8290;
  wire T8291;
  wire T8292;
  wire T8293;
  wire[46:0] T8294;
  wire[46:0] T8295;
  wire[46:0] T8296;
  wire[46:0] twiddle4_3_184_real;
  wire[46:0] T8297;
  wire[46:0] T8298;
  wire[46:0] T8299;
  wire[43:0] T8300;
  wire[43:0] T8301;
  wire[2:0] T8302;
  wire T8303;
  wire[46:0] twiddle4_3_185_real;
  wire[46:0] T8304;
  wire[46:0] T8305;
  wire[46:0] T8306;
  wire[44:0] T8307;
  wire[44:0] T8308;
  wire[1:0] T8309;
  wire T8310;
  wire T8311;
  wire[46:0] T8312;
  wire[46:0] twiddle4_3_186_real;
  wire[46:0] T8313;
  wire[46:0] T8314;
  wire[46:0] T8315;
  wire[44:0] T8316;
  wire[44:0] T8317;
  wire[1:0] T8318;
  wire T8319;
  wire[46:0] twiddle4_3_187_real;
  wire[46:0] T8320;
  wire[46:0] T8321;
  wire[46:0] T8322;
  wire[44:0] T8323;
  wire[44:0] T8324;
  wire[1:0] T8325;
  wire T8326;
  wire T8327;
  wire T8328;
  wire[46:0] T8329;
  wire[46:0] T8330;
  wire[46:0] twiddle4_3_188_real;
  wire[46:0] T8331;
  wire[46:0] T8332;
  wire[46:0] T8333;
  wire[44:0] T8334;
  wire[44:0] T8335;
  wire[1:0] T8336;
  wire T8337;
  wire[46:0] twiddle4_3_189_real;
  wire[46:0] T8338;
  wire[46:0] T8339;
  wire[46:0] T8340;
  wire[44:0] T8341;
  wire[44:0] T8342;
  wire[1:0] T8343;
  wire T8344;
  wire T8345;
  wire[46:0] T8346;
  wire[46:0] twiddle4_3_190_real;
  wire[46:0] T8347;
  wire[46:0] T8348;
  wire[46:0] T8349;
  wire[44:0] T8350;
  wire[44:0] T8351;
  wire[1:0] T8352;
  wire T8353;
  wire[46:0] twiddle4_3_191_real;
  wire[46:0] T8354;
  wire[46:0] T8355;
  wire[46:0] T8356;
  wire[44:0] T8357;
  wire[44:0] T8358;
  wire[1:0] T8359;
  wire T8360;
  wire T8361;
  wire T8362;
  wire T8363;
  wire T8364;
  wire T8365;
  wire T8366;
  wire[46:0] T8367;
  wire[46:0] T8368;
  wire[46:0] T8369;
  wire[46:0] T8370;
  wire[46:0] T8371;
  wire[46:0] T8372;
  wire[46:0] twiddle4_3_192_real;
  wire[46:0] T8373;
  wire[46:0] T8374;
  wire[46:0] T8375;
  wire[44:0] T8376;
  wire[44:0] T8377;
  wire[1:0] T8378;
  wire T8379;
  wire[46:0] twiddle4_3_193_real;
  wire[46:0] T8380;
  wire[46:0] T8381;
  wire[46:0] T8382;
  wire[44:0] T8383;
  wire[44:0] T8384;
  wire[1:0] T8385;
  wire T8386;
  wire T8387;
  wire[46:0] T8388;
  wire[46:0] twiddle4_3_194_real;
  wire[46:0] T8389;
  wire[46:0] T8390;
  wire[46:0] T8391;
  wire[44:0] T8392;
  wire[44:0] T8393;
  wire[1:0] T8394;
  wire T8395;
  wire[46:0] twiddle4_3_195_real;
  wire[46:0] T8396;
  wire[46:0] T8397;
  wire[46:0] T8398;
  wire[44:0] T8399;
  wire[44:0] T8400;
  wire[1:0] T8401;
  wire T8402;
  wire T8403;
  wire T8404;
  wire[46:0] T8405;
  wire[46:0] T8406;
  wire[46:0] twiddle4_3_196_real;
  wire[46:0] T8407;
  wire[46:0] T8408;
  wire[46:0] T8409;
  wire[44:0] T8410;
  wire[44:0] T8411;
  wire[1:0] T8412;
  wire T8413;
  wire[46:0] twiddle4_3_197_real;
  wire[46:0] T8414;
  wire[46:0] T8415;
  wire[46:0] T8416;
  wire[44:0] T8417;
  wire[44:0] T8418;
  wire[1:0] T8419;
  wire T8420;
  wire T8421;
  wire[46:0] T8422;
  wire[46:0] twiddle4_3_198_real;
  wire[46:0] T8423;
  wire[46:0] T8424;
  wire[46:0] T8425;
  wire[44:0] T8426;
  wire[44:0] T8427;
  wire[1:0] T8428;
  wire T8429;
  wire[46:0] twiddle4_3_199_real;
  wire[46:0] T8430;
  wire[46:0] T8431;
  wire[46:0] T8432;
  wire[45:0] T8433;
  wire[45:0] T8434;
  wire T8435;
  wire T8436;
  wire T8437;
  wire T8438;
  wire[46:0] T8439;
  wire[46:0] T8440;
  wire[46:0] T8441;
  wire[46:0] twiddle4_3_200_real;
  wire[46:0] T8442;
  wire[46:0] T8443;
  wire[46:0] T8444;
  wire[45:0] T8445;
  wire[45:0] T8446;
  wire T8447;
  wire[46:0] twiddle4_3_201_real;
  wire[46:0] T8448;
  wire[46:0] T8449;
  wire[46:0] T8450;
  wire[45:0] T8451;
  wire[45:0] T8452;
  wire T8453;
  wire T8454;
  wire[46:0] T8455;
  wire[46:0] twiddle4_3_202_real;
  wire[46:0] T8456;
  wire[46:0] T8457;
  wire[46:0] T8458;
  wire[45:0] T8459;
  wire[45:0] T8460;
  wire T8461;
  wire[46:0] twiddle4_3_203_real;
  wire[46:0] T8462;
  wire[46:0] T8463;
  wire[46:0] T8464;
  wire[45:0] T8465;
  wire[45:0] T8466;
  wire T8467;
  wire T8468;
  wire T8469;
  wire[46:0] T8470;
  wire[46:0] T8471;
  wire[46:0] twiddle4_3_204_real;
  wire[46:0] T8472;
  wire[46:0] T8473;
  wire[46:0] T8474;
  wire[45:0] T8475;
  wire[45:0] T8476;
  wire T8477;
  wire[46:0] twiddle4_3_205_real;
  wire[46:0] T8478;
  wire[46:0] T8479;
  wire[46:0] T8480;
  wire[45:0] T8481;
  wire[45:0] T8482;
  wire T8483;
  wire T8484;
  wire[46:0] T8485;
  wire[46:0] twiddle4_3_206_real;
  wire[46:0] T8486;
  wire[46:0] T8487;
  wire[46:0] T8488;
  wire[45:0] T8489;
  wire[45:0] T8490;
  wire T8491;
  wire[46:0] twiddle4_3_207_real;
  wire[46:0] T8492;
  wire[46:0] T8493;
  wire[46:0] T8494;
  wire[45:0] T8495;
  wire[45:0] T8496;
  wire T8497;
  wire T8498;
  wire T8499;
  wire T8500;
  wire T8501;
  wire[46:0] T8502;
  wire[46:0] T8503;
  wire[46:0] T8504;
  wire[46:0] T8505;
  wire[46:0] twiddle4_3_208_real;
  wire[46:0] T8506;
  wire[46:0] T8507;
  wire[46:0] T8508;
  wire[45:0] T8509;
  wire[45:0] T8510;
  wire T8511;
  wire[46:0] twiddle4_3_209_real;
  wire[46:0] T8512;
  wire[46:0] T8513;
  wire[46:0] T8514;
  wire[45:0] T8515;
  wire[45:0] T8516;
  wire T8517;
  wire T8518;
  wire[46:0] T8519;
  wire[46:0] twiddle4_3_210_real;
  wire[46:0] T8520;
  wire[46:0] T8521;
  wire[46:0] T8522;
  wire[45:0] T8523;
  wire[45:0] T8524;
  wire T8525;
  wire[46:0] twiddle4_3_211_real;
  wire[46:0] T8526;
  wire[46:0] T8527;
  wire[46:0] T8528;
  wire[45:0] T8529;
  wire[45:0] T8530;
  wire T8531;
  wire T8532;
  wire T8533;
  wire[46:0] T8534;
  wire[46:0] T8535;
  wire[46:0] twiddle4_3_212_real;
  wire[46:0] T8536;
  wire[46:0] T8537;
  wire[46:0] T8538;
  wire[45:0] T8539;
  wire[45:0] T8540;
  wire T8541;
  wire[46:0] twiddle4_3_213_real;
  wire[46:0] T8542;
  wire[46:0] T8543;
  wire[46:0] T8544;
  wire[45:0] T8545;
  wire[45:0] T8546;
  wire T8547;
  wire T8548;
  wire[46:0] T8549;
  wire[46:0] twiddle4_3_214_real;
  wire[46:0] T8550;
  wire[46:0] T8551;
  wire[46:0] T8552;
  wire[45:0] T8553;
  wire[45:0] T8554;
  wire T8555;
  wire[46:0] twiddle4_3_215_real;
  wire[46:0] T8556;
  wire[46:0] T8557;
  wire[46:0] T8558;
  wire[45:0] T8559;
  wire[45:0] T8560;
  wire T8561;
  wire T8562;
  wire T8563;
  wire T8564;
  wire[46:0] T8565;
  wire[46:0] T8566;
  wire[46:0] T8567;
  wire[46:0] twiddle4_3_216_real;
  wire[46:0] T8568;
  wire[46:0] T8569;
  wire[46:0] T8570;
  wire[45:0] T8571;
  wire[45:0] T8572;
  wire T8573;
  wire[46:0] twiddle4_3_217_real;
  wire[46:0] T8574;
  wire[46:0] T8575;
  wire[46:0] T8576;
  wire[45:0] T8577;
  wire[45:0] T8578;
  wire T8579;
  wire T8580;
  wire[46:0] T8581;
  wire[46:0] twiddle4_3_218_real;
  wire[46:0] T8582;
  wire[46:0] T8583;
  wire[46:0] T8584;
  wire[45:0] T8585;
  wire[45:0] T8586;
  wire T8587;
  wire[46:0] twiddle4_3_219_real;
  wire[46:0] T8588;
  wire[46:0] T8589;
  wire[46:0] T8590;
  wire[45:0] T8591;
  wire[45:0] T8592;
  wire T8593;
  wire T8594;
  wire T8595;
  wire[46:0] T8596;
  wire[46:0] T8597;
  wire[46:0] twiddle4_3_220_real;
  wire[46:0] T8598;
  wire[46:0] T8599;
  wire[46:0] T8600;
  wire[45:0] T8601;
  wire[45:0] T8602;
  wire T8603;
  wire[46:0] twiddle4_3_221_real;
  wire[46:0] T8604;
  wire[46:0] T8605;
  wire[46:0] T8606;
  wire[45:0] T8607;
  wire[45:0] T8608;
  wire T8609;
  wire T8610;
  wire[46:0] T8611;
  wire[46:0] twiddle4_3_222_real;
  wire[46:0] T8612;
  wire[46:0] T8613;
  wire[46:0] T8614;
  wire[45:0] T8615;
  wire[45:0] T8616;
  wire T8617;
  wire[46:0] twiddle4_3_223_real;
  wire[46:0] T8618;
  wire[46:0] T8619;
  wire[46:0] T8620;
  wire[45:0] T8621;
  wire[45:0] T8622;
  wire T8623;
  wire T8624;
  wire T8625;
  wire T8626;
  wire T8627;
  wire T8628;
  wire[46:0] T8629;
  wire[46:0] T8630;
  wire[46:0] T8631;
  wire[46:0] T8632;
  wire[46:0] T8633;
  wire[46:0] twiddle4_3_224_real;
  wire[46:0] T8634;
  wire[46:0] T8635;
  wire[46:0] T8636;
  wire[45:0] T8637;
  wire[45:0] T8638;
  wire T8639;
  wire[46:0] twiddle4_3_225_real;
  wire[46:0] T8640;
  wire[46:0] T8641;
  wire[46:0] T8642;
  wire[45:0] T8643;
  wire[45:0] T8644;
  wire T8645;
  wire T8646;
  wire[46:0] T8647;
  wire[46:0] twiddle4_3_226_real;
  wire[46:0] T8648;
  wire[46:0] T8649;
  wire[46:0] T8650;
  wire[45:0] T8651;
  wire[45:0] T8652;
  wire T8653;
  wire[46:0] twiddle4_3_227_real;
  wire[46:0] T8654;
  wire[46:0] T8655;
  wire[46:0] T8656;
  wire[45:0] T8657;
  wire[45:0] T8658;
  wire T8659;
  wire T8660;
  wire T8661;
  wire[46:0] T8662;
  wire[46:0] T8663;
  wire[46:0] twiddle4_3_228_real;
  wire[46:0] T8664;
  wire[46:0] T8665;
  wire[46:0] T8666;
  wire[46:0] T8667;
  wire[46:0] twiddle4_3_229_real;
  wire[46:0] T8668;
  wire[46:0] T8669;
  wire[46:0] T8670;
  wire[46:0] T8671;
  wire T8672;
  wire[46:0] T8673;
  wire[46:0] twiddle4_3_230_real;
  wire[46:0] T8674;
  wire[46:0] T8675;
  wire[46:0] T8676;
  wire[46:0] T8677;
  wire[46:0] twiddle4_3_231_real;
  wire[46:0] T8678;
  wire[46:0] T8679;
  wire[46:0] T8680;
  wire[46:0] T8681;
  wire T8682;
  wire T8683;
  wire T8684;
  wire[46:0] T8685;
  wire[46:0] T8686;
  wire[46:0] T8687;
  wire[46:0] twiddle4_3_232_real;
  wire[46:0] T8688;
  wire[46:0] T8689;
  wire[46:0] T8690;
  wire[46:0] T8691;
  wire[46:0] twiddle4_3_233_real;
  wire[46:0] T8692;
  wire[46:0] T8693;
  wire[46:0] T8694;
  wire[46:0] T8695;
  wire T8696;
  wire[46:0] T8697;
  wire[46:0] twiddle4_3_234_real;
  wire[46:0] T8698;
  wire[46:0] T8699;
  wire[46:0] T8700;
  wire[46:0] T8701;
  wire[46:0] twiddle4_3_235_real;
  wire[46:0] T8702;
  wire[46:0] T8703;
  wire[46:0] T8704;
  wire[46:0] T8705;
  wire T8706;
  wire T8707;
  wire[46:0] T8708;
  wire[46:0] T8709;
  wire[46:0] twiddle4_3_236_real;
  wire[46:0] T8710;
  wire[46:0] T8711;
  wire[46:0] T8712;
  wire[46:0] T8713;
  wire[46:0] twiddle4_3_237_real;
  wire[46:0] T8714;
  wire[46:0] T8715;
  wire[46:0] T8716;
  wire[46:0] T8717;
  wire T8718;
  wire[46:0] T8719;
  wire[46:0] twiddle4_3_238_real;
  wire[46:0] T8720;
  wire[46:0] T8721;
  wire[46:0] T8722;
  wire[46:0] T8723;
  wire[46:0] twiddle4_3_239_real;
  wire[46:0] T8724;
  wire[46:0] T8725;
  wire[46:0] T8726;
  wire[46:0] T8727;
  wire T8728;
  wire T8729;
  wire T8730;
  wire T8731;
  wire[46:0] T8732;
  wire[46:0] T8733;
  wire[46:0] T8734;
  wire[46:0] T8735;
  wire[46:0] twiddle4_3_240_real;
  wire[46:0] T8736;
  wire[46:0] T8737;
  wire[46:0] T8738;
  wire[46:0] T8739;
  wire[46:0] twiddle4_3_241_real;
  wire[46:0] T8740;
  wire[46:0] T8741;
  wire[46:0] T8742;
  wire[46:0] T8743;
  wire T8744;
  wire[46:0] T8745;
  wire[46:0] twiddle4_3_242_real;
  wire[46:0] T8746;
  wire[46:0] T8747;
  wire[46:0] T8748;
  wire[46:0] T8749;
  wire[46:0] twiddle4_3_243_real;
  wire[46:0] T8750;
  wire[46:0] T8751;
  wire[46:0] T8752;
  wire[46:0] T8753;
  wire T8754;
  wire T8755;
  wire[46:0] T8756;
  wire[46:0] T8757;
  wire[46:0] twiddle4_3_244_real;
  wire[46:0] T8758;
  wire[46:0] T8759;
  wire[46:0] T8760;
  wire[46:0] T8761;
  wire[46:0] twiddle4_3_245_real;
  wire[46:0] T8762;
  wire[46:0] T8763;
  wire[46:0] T8764;
  wire[46:0] T8765;
  wire T8766;
  wire[46:0] T8767;
  wire[46:0] twiddle4_3_246_real;
  wire[46:0] T8768;
  wire[46:0] T8769;
  wire[46:0] T8770;
  wire[46:0] T8771;
  wire[46:0] twiddle4_3_247_real;
  wire[46:0] T8772;
  wire[46:0] T8773;
  wire[46:0] T8774;
  wire[46:0] T8775;
  wire T8776;
  wire T8777;
  wire T8778;
  wire[46:0] T8779;
  wire[46:0] T8780;
  wire[46:0] T8781;
  wire[46:0] twiddle4_3_248_real;
  wire[46:0] T8782;
  wire[46:0] T8783;
  wire[46:0] T8784;
  wire[46:0] T8785;
  wire[46:0] twiddle4_3_249_real;
  wire[46:0] T8786;
  wire[46:0] T8787;
  wire[46:0] T8788;
  wire[46:0] T8789;
  wire T8790;
  wire[46:0] T8791;
  wire[46:0] twiddle4_3_250_real;
  wire[46:0] T8792;
  wire[46:0] T8793;
  wire[46:0] T8794;
  wire[46:0] T8795;
  wire[46:0] twiddle4_3_251_real;
  wire[46:0] T8796;
  wire[46:0] T8797;
  wire[46:0] T8798;
  wire[46:0] T8799;
  wire T8800;
  wire T8801;
  wire[46:0] T8802;
  wire[46:0] T8803;
  wire[46:0] twiddle4_3_252_real;
  wire[46:0] T8804;
  wire[46:0] T8805;
  wire[46:0] T8806;
  wire[46:0] T8807;
  wire[46:0] twiddle4_3_253_real;
  wire[46:0] T8808;
  wire[46:0] T8809;
  wire[46:0] T8810;
  wire[46:0] T8811;
  wire T8812;
  wire[46:0] T8813;
  wire[46:0] twiddle4_3_254_real;
  wire[46:0] T8814;
  wire[46:0] T8815;
  wire[46:0] T8816;
  wire[46:0] T8817;
  wire[46:0] twiddle4_3_255_real;
  wire[46:0] T8818;
  wire[46:0] T8819;
  wire[46:0] T8820;
  wire[46:0] T8821;
  wire T8822;
  wire T8823;
  wire T8824;
  wire T8825;
  wire T8826;
  wire T8827;
  wire T8828;
  wire T8829;
  wire T8830;
  wire[47:0] T8831;
  wire[46:0] T8832;
  wire[46:0] T8833;
  wire[46:0] T8834;
  wire[46:0] T8835;
  wire[46:0] T8836;
  wire[46:0] T8837;
  wire[46:0] T8838;
  wire[46:0] T8839;
  wire[46:0] twiddle4_3_256_real;
  wire[46:0] T8840;
  wire[46:0] T8841;
  wire[46:0] T8842;
  wire[46:0] T8843;
  wire[46:0] twiddle4_3_257_real;
  wire[46:0] T8844;
  wire[46:0] T8845;
  wire[46:0] T8846;
  wire[46:0] T8847;
  wire T8848;
  wire[46:0] T8849;
  wire[46:0] twiddle4_3_258_real;
  wire[46:0] T8850;
  wire[46:0] T8851;
  wire[46:0] T8852;
  wire[46:0] T8853;
  wire[46:0] twiddle4_3_259_real;
  wire[46:0] T8854;
  wire[46:0] T8855;
  wire[46:0] T8856;
  wire[46:0] T8857;
  wire T8858;
  wire T8859;
  wire[46:0] T8860;
  wire[46:0] T8861;
  wire[46:0] twiddle4_3_260_real;
  wire[46:0] T8862;
  wire[46:0] T8863;
  wire[46:0] T8864;
  wire[46:0] T8865;
  wire[46:0] twiddle4_3_261_real;
  wire[46:0] T8866;
  wire[46:0] T8867;
  wire[46:0] T8868;
  wire[46:0] T8869;
  wire T8870;
  wire[46:0] T8871;
  wire[46:0] twiddle4_3_262_real;
  wire[46:0] T8872;
  wire[46:0] T8873;
  wire[46:0] T8874;
  wire[46:0] T8875;
  wire[46:0] twiddle4_3_263_real;
  wire[46:0] T8876;
  wire[46:0] T8877;
  wire[46:0] T8878;
  wire[46:0] T8879;
  wire T8880;
  wire T8881;
  wire T8882;
  wire[46:0] T8883;
  wire[46:0] T8884;
  wire[46:0] T8885;
  wire[46:0] twiddle4_3_264_real;
  wire[46:0] T8886;
  wire[46:0] T8887;
  wire[46:0] T8888;
  wire[46:0] T8889;
  wire[46:0] twiddle4_3_265_real;
  wire[46:0] T8890;
  wire[46:0] T8891;
  wire[46:0] T8892;
  wire[46:0] T8893;
  wire T8894;
  wire[46:0] T8895;
  wire[46:0] twiddle4_3_266_real;
  wire[46:0] T8896;
  wire[46:0] T8897;
  wire[46:0] T8898;
  wire[46:0] T8899;
  wire[46:0] twiddle4_3_267_real;
  wire[46:0] T8900;
  wire[46:0] T8901;
  wire[46:0] T8902;
  wire[46:0] T8903;
  wire T8904;
  wire T8905;
  wire[46:0] T8906;
  wire[46:0] T8907;
  wire[46:0] twiddle4_3_268_real;
  wire[46:0] T8908;
  wire[46:0] T8909;
  wire[46:0] T8910;
  wire[46:0] T8911;
  wire[46:0] twiddle4_3_269_real;
  wire[46:0] T8912;
  wire[46:0] T8913;
  wire[46:0] T8914;
  wire[46:0] T8915;
  wire T8916;
  wire[46:0] T8917;
  wire[46:0] twiddle4_3_270_real;
  wire[46:0] T8918;
  wire[46:0] T8919;
  wire[46:0] T8920;
  wire[46:0] T8921;
  wire[46:0] twiddle4_3_271_real;
  wire[46:0] T8922;
  wire[46:0] T8923;
  wire[46:0] T8924;
  wire[46:0] T8925;
  wire T8926;
  wire T8927;
  wire T8928;
  wire T8929;
  wire[46:0] T8930;
  wire[46:0] T8931;
  wire[46:0] T8932;
  wire[46:0] T8933;
  wire[46:0] twiddle4_3_272_real;
  wire[46:0] T8934;
  wire[46:0] T8935;
  wire[46:0] T8936;
  wire[46:0] T8937;
  wire[46:0] twiddle4_3_273_real;
  wire[46:0] T8938;
  wire[46:0] T8939;
  wire[46:0] T8940;
  wire[46:0] T8941;
  wire T8942;
  wire[46:0] T8943;
  wire[46:0] twiddle4_3_274_real;
  wire[46:0] T8944;
  wire[46:0] T8945;
  wire[46:0] T8946;
  wire[46:0] T8947;
  wire[46:0] twiddle4_3_275_real;
  wire[46:0] T8948;
  wire[46:0] T8949;
  wire[46:0] T8950;
  wire[46:0] T8951;
  wire T8952;
  wire T8953;
  wire[46:0] T8954;
  wire[46:0] T8955;
  wire[46:0] twiddle4_3_276_real;
  wire[46:0] T8956;
  wire[46:0] T8957;
  wire[46:0] T8958;
  wire[46:0] T8959;
  wire[46:0] twiddle4_3_277_real;
  wire[46:0] T8960;
  wire[46:0] T8961;
  wire[46:0] T8962;
  wire[46:0] T8963;
  wire T8964;
  wire[46:0] T8965;
  wire[46:0] twiddle4_3_278_real;
  wire[46:0] T8966;
  wire[46:0] T8967;
  wire[46:0] T8968;
  wire[46:0] T8969;
  wire[46:0] twiddle4_3_279_real;
  wire[46:0] T8970;
  wire[46:0] T8971;
  wire[46:0] T8972;
  wire[46:0] T8973;
  wire T8974;
  wire T8975;
  wire T8976;
  wire[46:0] T8977;
  wire[46:0] T8978;
  wire[46:0] T8979;
  wire[46:0] twiddle4_3_280_real;
  wire[46:0] T8980;
  wire[46:0] T8981;
  wire[46:0] T8982;
  wire[46:0] T8983;
  wire[46:0] twiddle4_3_281_real;
  wire[46:0] T8984;
  wire[46:0] T8985;
  wire[46:0] T8986;
  wire[46:0] T8987;
  wire T8988;
  wire[46:0] T8989;
  wire[46:0] twiddle4_3_282_real;
  wire[46:0] T8990;
  wire[46:0] T8991;
  wire[46:0] T8992;
  wire[46:0] T8993;
  wire[46:0] twiddle4_3_283_real;
  wire[46:0] T8994;
  wire[46:0] T8995;
  wire[46:0] T8996;
  wire[46:0] T8997;
  wire T8998;
  wire T8999;
  wire[46:0] T9000;
  wire[46:0] T9001;
  wire[46:0] twiddle4_3_284_real;
  wire[46:0] T9002;
  wire[46:0] T9003;
  wire[46:0] T9004;
  wire[46:0] T9005;
  wire[46:0] twiddle4_3_285_real;
  wire[46:0] T9006;
  wire[45:0] T9007;
  wire[45:0] T9008;
  wire T9009;
  wire[46:0] T9010;
  wire[46:0] T9011;
  wire T9012;
  wire[46:0] T9013;
  wire[46:0] twiddle4_3_286_real;
  wire[46:0] T9014;
  wire[45:0] T9015;
  wire[45:0] T9016;
  wire T9017;
  wire[46:0] T9018;
  wire[46:0] T9019;
  wire[46:0] twiddle4_3_287_real;
  wire[46:0] T9020;
  wire[45:0] T9021;
  wire[45:0] T9022;
  wire T9023;
  wire[46:0] T9024;
  wire[46:0] T9025;
  wire T9026;
  wire T9027;
  wire T9028;
  wire T9029;
  wire T9030;
  wire[46:0] T9031;
  wire[46:0] T9032;
  wire[46:0] T9033;
  wire[46:0] T9034;
  wire[46:0] T9035;
  wire[46:0] twiddle4_3_288_real;
  wire[46:0] T9036;
  wire[45:0] T9037;
  wire[45:0] T9038;
  wire T9039;
  wire[46:0] T9040;
  wire[46:0] T9041;
  wire[46:0] twiddle4_3_289_real;
  wire[46:0] T9042;
  wire[45:0] T9043;
  wire[45:0] T9044;
  wire T9045;
  wire[46:0] T9046;
  wire[46:0] T9047;
  wire T9048;
  wire[46:0] T9049;
  wire[46:0] twiddle4_3_290_real;
  wire[46:0] T9050;
  wire[45:0] T9051;
  wire[45:0] T9052;
  wire T9053;
  wire[46:0] T9054;
  wire[46:0] T9055;
  wire[46:0] twiddle4_3_291_real;
  wire[46:0] T9056;
  wire[45:0] T9057;
  wire[45:0] T9058;
  wire T9059;
  wire[46:0] T9060;
  wire[46:0] T9061;
  wire T9062;
  wire T9063;
  wire[46:0] T9064;
  wire[46:0] T9065;
  wire[46:0] twiddle4_3_292_real;
  wire[46:0] T9066;
  wire[45:0] T9067;
  wire[45:0] T9068;
  wire T9069;
  wire[46:0] T9070;
  wire[46:0] T9071;
  wire[46:0] twiddle4_3_293_real;
  wire[46:0] T9072;
  wire[45:0] T9073;
  wire[45:0] T9074;
  wire T9075;
  wire[46:0] T9076;
  wire[46:0] T9077;
  wire T9078;
  wire[46:0] T9079;
  wire[46:0] twiddle4_3_294_real;
  wire[46:0] T9080;
  wire[45:0] T9081;
  wire[45:0] T9082;
  wire T9083;
  wire[46:0] T9084;
  wire[46:0] T9085;
  wire[46:0] twiddle4_3_295_real;
  wire[46:0] T9086;
  wire[45:0] T9087;
  wire[45:0] T9088;
  wire T9089;
  wire[46:0] T9090;
  wire[46:0] T9091;
  wire T9092;
  wire T9093;
  wire T9094;
  wire[46:0] T9095;
  wire[46:0] T9096;
  wire[46:0] T9097;
  wire[46:0] twiddle4_3_296_real;
  wire[46:0] T9098;
  wire[45:0] T9099;
  wire[45:0] T9100;
  wire T9101;
  wire[46:0] T9102;
  wire[46:0] T9103;
  wire[46:0] twiddle4_3_297_real;
  wire[46:0] T9104;
  wire[45:0] T9105;
  wire[45:0] T9106;
  wire T9107;
  wire[46:0] T9108;
  wire[46:0] T9109;
  wire T9110;
  wire[46:0] T9111;
  wire[46:0] twiddle4_3_298_real;
  wire[46:0] T9112;
  wire[45:0] T9113;
  wire[45:0] T9114;
  wire T9115;
  wire[46:0] T9116;
  wire[46:0] T9117;
  wire[46:0] twiddle4_3_299_real;
  wire[46:0] T9118;
  wire[45:0] T9119;
  wire[45:0] T9120;
  wire T9121;
  wire[46:0] T9122;
  wire[46:0] T9123;
  wire T9124;
  wire T9125;
  wire[46:0] T9126;
  wire[46:0] T9127;
  wire[46:0] twiddle4_3_300_real;
  wire[46:0] T9128;
  wire[45:0] T9129;
  wire[45:0] T9130;
  wire T9131;
  wire[46:0] T9132;
  wire[46:0] T9133;
  wire[46:0] twiddle4_3_301_real;
  wire[46:0] T9134;
  wire[45:0] T9135;
  wire[45:0] T9136;
  wire T9137;
  wire[46:0] T9138;
  wire[46:0] T9139;
  wire T9140;
  wire[46:0] T9141;
  wire[46:0] twiddle4_3_302_real;
  wire[46:0] T9142;
  wire[45:0] T9143;
  wire[45:0] T9144;
  wire T9145;
  wire[46:0] T9146;
  wire[46:0] T9147;
  wire[46:0] twiddle4_3_303_real;
  wire[46:0] T9148;
  wire[45:0] T9149;
  wire[45:0] T9150;
  wire T9151;
  wire[46:0] T9152;
  wire[46:0] T9153;
  wire T9154;
  wire T9155;
  wire T9156;
  wire T9157;
  wire[46:0] T9158;
  wire[46:0] T9159;
  wire[46:0] T9160;
  wire[46:0] T9161;
  wire[46:0] twiddle4_3_304_real;
  wire[46:0] T9162;
  wire[45:0] T9163;
  wire[45:0] T9164;
  wire T9165;
  wire[46:0] T9166;
  wire[46:0] T9167;
  wire[46:0] twiddle4_3_305_real;
  wire[46:0] T9168;
  wire[45:0] T9169;
  wire[45:0] T9170;
  wire T9171;
  wire[46:0] T9172;
  wire[46:0] T9173;
  wire T9174;
  wire[46:0] T9175;
  wire[46:0] twiddle4_3_306_real;
  wire[46:0] T9176;
  wire[45:0] T9177;
  wire[45:0] T9178;
  wire T9179;
  wire[46:0] T9180;
  wire[46:0] T9181;
  wire[46:0] twiddle4_3_307_real;
  wire[46:0] T9182;
  wire[45:0] T9183;
  wire[45:0] T9184;
  wire T9185;
  wire[46:0] T9186;
  wire[46:0] T9187;
  wire T9188;
  wire T9189;
  wire[46:0] T9190;
  wire[46:0] T9191;
  wire[46:0] twiddle4_3_308_real;
  wire[46:0] T9192;
  wire[45:0] T9193;
  wire[45:0] T9194;
  wire T9195;
  wire[46:0] T9196;
  wire[46:0] T9197;
  wire[46:0] twiddle4_3_309_real;
  wire[46:0] T9198;
  wire[45:0] T9199;
  wire[45:0] T9200;
  wire T9201;
  wire[46:0] T9202;
  wire[46:0] T9203;
  wire T9204;
  wire[46:0] T9205;
  wire[46:0] twiddle4_3_310_real;
  wire[46:0] T9206;
  wire[45:0] T9207;
  wire[45:0] T9208;
  wire T9209;
  wire[46:0] T9210;
  wire[46:0] T9211;
  wire[46:0] twiddle4_3_311_real;
  wire[46:0] T9212;
  wire[45:0] T9213;
  wire[45:0] T9214;
  wire T9215;
  wire[46:0] T9216;
  wire[46:0] T9217;
  wire T9218;
  wire T9219;
  wire T9220;
  wire[46:0] T9221;
  wire[46:0] T9222;
  wire[46:0] T9223;
  wire[46:0] twiddle4_3_312_real;
  wire[46:0] T9224;
  wire[45:0] T9225;
  wire[45:0] T9226;
  wire T9227;
  wire[46:0] T9228;
  wire[46:0] T9229;
  wire[46:0] twiddle4_3_313_real;
  wire[46:0] T9230;
  wire[45:0] T9231;
  wire[45:0] T9232;
  wire T9233;
  wire[46:0] T9234;
  wire[46:0] T9235;
  wire T9236;
  wire[46:0] T9237;
  wire[46:0] twiddle4_3_314_real;
  wire[46:0] T9238;
  wire[44:0] T9239;
  wire[44:0] T9240;
  wire[1:0] T9241;
  wire T9242;
  wire[46:0] T9243;
  wire[46:0] T9244;
  wire[46:0] twiddle4_3_315_real;
  wire[46:0] T9245;
  wire[44:0] T9246;
  wire[44:0] T9247;
  wire[1:0] T9248;
  wire T9249;
  wire[46:0] T9250;
  wire[46:0] T9251;
  wire T9252;
  wire T9253;
  wire[46:0] T9254;
  wire[46:0] T9255;
  wire[46:0] twiddle4_3_316_real;
  wire[46:0] T9256;
  wire[44:0] T9257;
  wire[44:0] T9258;
  wire[1:0] T9259;
  wire T9260;
  wire[46:0] T9261;
  wire[46:0] T9262;
  wire[46:0] twiddle4_3_317_real;
  wire[46:0] T9263;
  wire[44:0] T9264;
  wire[44:0] T9265;
  wire[1:0] T9266;
  wire T9267;
  wire[46:0] T9268;
  wire[46:0] T9269;
  wire T9270;
  wire[46:0] T9271;
  wire[46:0] twiddle4_3_318_real;
  wire[46:0] T9272;
  wire[44:0] T9273;
  wire[44:0] T9274;
  wire[1:0] T9275;
  wire T9276;
  wire[46:0] T9277;
  wire[46:0] T9278;
  wire[46:0] twiddle4_3_319_real;
  wire[46:0] T9279;
  wire[44:0] T9280;
  wire[44:0] T9281;
  wire[1:0] T9282;
  wire T9283;
  wire[46:0] T9284;
  wire[46:0] T9285;
  wire T9286;
  wire T9287;
  wire T9288;
  wire T9289;
  wire T9290;
  wire T9291;
  wire[46:0] T9292;
  wire[46:0] T9293;
  wire[46:0] T9294;
  wire[46:0] T9295;
  wire[46:0] T9296;
  wire[46:0] T9297;
  wire[46:0] twiddle4_3_320_real;
  wire[46:0] T9298;
  wire[44:0] T9299;
  wire[44:0] T9300;
  wire[1:0] T9301;
  wire T9302;
  wire[46:0] T9303;
  wire[46:0] T9304;
  wire[46:0] twiddle4_3_321_real;
  wire[46:0] T9305;
  wire[44:0] T9306;
  wire[44:0] T9307;
  wire[1:0] T9308;
  wire T9309;
  wire[46:0] T9310;
  wire[46:0] T9311;
  wire T9312;
  wire[46:0] T9313;
  wire[46:0] twiddle4_3_322_real;
  wire[46:0] T9314;
  wire[44:0] T9315;
  wire[44:0] T9316;
  wire[1:0] T9317;
  wire T9318;
  wire[46:0] T9319;
  wire[46:0] T9320;
  wire[46:0] twiddle4_3_323_real;
  wire[46:0] T9321;
  wire[44:0] T9322;
  wire[44:0] T9323;
  wire[1:0] T9324;
  wire T9325;
  wire[46:0] T9326;
  wire[46:0] T9327;
  wire T9328;
  wire T9329;
  wire[46:0] T9330;
  wire[46:0] T9331;
  wire[46:0] twiddle4_3_324_real;
  wire[46:0] T9332;
  wire[44:0] T9333;
  wire[44:0] T9334;
  wire[1:0] T9335;
  wire T9336;
  wire[46:0] T9337;
  wire[46:0] T9338;
  wire[46:0] twiddle4_3_325_real;
  wire[46:0] T9339;
  wire[44:0] T9340;
  wire[44:0] T9341;
  wire[1:0] T9342;
  wire T9343;
  wire[46:0] T9344;
  wire[46:0] T9345;
  wire T9346;
  wire[46:0] T9347;
  wire[46:0] twiddle4_3_326_real;
  wire[46:0] T9348;
  wire[44:0] T9349;
  wire[44:0] T9350;
  wire[1:0] T9351;
  wire T9352;
  wire[46:0] T9353;
  wire[46:0] T9354;
  wire[46:0] twiddle4_3_327_real;
  wire[46:0] T9355;
  wire[44:0] T9356;
  wire[44:0] T9357;
  wire[1:0] T9358;
  wire T9359;
  wire[46:0] T9360;
  wire[46:0] T9361;
  wire T9362;
  wire T9363;
  wire T9364;
  wire[46:0] T9365;
  wire[46:0] T9366;
  wire[46:0] T9367;
  wire[46:0] twiddle4_3_328_real;
  wire[46:0] T9368;
  wire[43:0] T9369;
  wire[43:0] T9370;
  wire[2:0] T9371;
  wire T9372;
  wire[46:0] T9373;
  wire[46:0] T9374;
  wire[46:0] twiddle4_3_329_real;
  wire[46:0] T9375;
  wire[43:0] T9376;
  wire[43:0] T9377;
  wire[2:0] T9378;
  wire T9379;
  wire[46:0] T9380;
  wire[46:0] T9381;
  wire T9382;
  wire[46:0] T9383;
  wire[46:0] twiddle4_3_330_real;
  wire[46:0] T9384;
  wire[43:0] T9385;
  wire[43:0] T9386;
  wire[2:0] T9387;
  wire T9388;
  wire[46:0] T9389;
  wire[46:0] T9390;
  wire[46:0] twiddle4_3_331_real;
  wire[46:0] T9391;
  wire[43:0] T9392;
  wire[43:0] T9393;
  wire[2:0] T9394;
  wire T9395;
  wire[46:0] T9396;
  wire[46:0] T9397;
  wire T9398;
  wire T9399;
  wire[46:0] T9400;
  wire[46:0] T9401;
  wire[46:0] twiddle4_3_332_real;
  wire[46:0] T9402;
  wire[43:0] T9403;
  wire[43:0] T9404;
  wire[2:0] T9405;
  wire T9406;
  wire[46:0] T9407;
  wire[46:0] T9408;
  wire[46:0] twiddle4_3_333_real;
  wire[46:0] T9409;
  wire[43:0] T9410;
  wire[43:0] T9411;
  wire[2:0] T9412;
  wire T9413;
  wire[46:0] T9414;
  wire[46:0] T9415;
  wire T9416;
  wire[46:0] T9417;
  wire[46:0] twiddle4_3_334_real;
  wire[46:0] T9418;
  wire[43:0] T9419;
  wire[43:0] T9420;
  wire[2:0] T9421;
  wire T9422;
  wire[46:0] T9423;
  wire[46:0] T9424;
  wire[46:0] twiddle4_3_335_real;
  wire[46:0] T9425;
  wire[42:0] T9426;
  wire[42:0] T9427;
  wire[3:0] T9428;
  wire T9429;
  wire[46:0] T9430;
  wire[46:0] T9431;
  wire T9432;
  wire T9433;
  wire T9434;
  wire T9435;
  wire[46:0] T9436;
  wire[46:0] T9437;
  wire[46:0] T9438;
  wire[46:0] T9439;
  wire[46:0] twiddle4_3_336_real;
  wire[46:0] T9440;
  wire[42:0] T9441;
  wire[42:0] T9442;
  wire[3:0] T9443;
  wire T9444;
  wire[46:0] T9445;
  wire[46:0] T9446;
  wire[46:0] twiddle4_3_337_real;
  wire[46:0] T9447;
  wire[42:0] T9448;
  wire[42:0] T9449;
  wire[3:0] T9450;
  wire T9451;
  wire[46:0] T9452;
  wire[46:0] T9453;
  wire T9454;
  wire[46:0] T9455;
  wire[46:0] twiddle4_3_338_real;
  wire[46:0] T9456;
  wire[41:0] T9457;
  wire[41:0] T9458;
  wire[4:0] T9459;
  wire T9460;
  wire[46:0] T9461;
  wire[46:0] T9462;
  wire[46:0] twiddle4_3_339_real;
  wire[46:0] T9463;
  wire[41:0] T9464;
  wire[41:0] T9465;
  wire[4:0] T9466;
  wire T9467;
  wire[46:0] T9468;
  wire[46:0] T9469;
  wire T9470;
  wire T9471;
  wire[46:0] T9472;
  wire[46:0] T9473;
  wire[46:0] twiddle4_3_340_real;
  wire[46:0] T9474;
  wire[40:0] T9475;
  wire[40:0] T9476;
  wire[5:0] T9477;
  wire T9478;
  wire[46:0] T9479;
  wire[46:0] T9480;
  wire[46:0] twiddle4_3_341_real;
  wire[46:0] T9481;
  wire[38:0] T9482;
  wire[38:0] T9483;
  wire[7:0] T9484;
  wire T9485;
  wire[46:0] T9486;
  wire[46:0] T9487;
  wire T9488;
  wire[46:0] T9489;
  wire[46:0] twiddle4_3_342_real;
  wire[46:0] T9490;
  wire[39:0] T9491;
  wire[39:0] T9492;
  wire[6:0] T9493;
  wire T9494;
  wire[46:0] T9495;
  wire[46:0] T9496;
  wire[46:0] twiddle4_3_343_real;
  wire[46:0] T9497;
  wire[40:0] T9498;
  wire[40:0] T9499;
  wire[5:0] T9500;
  wire T9501;
  wire[46:0] T9502;
  wire[46:0] T9503;
  wire T9504;
  wire T9505;
  wire T9506;
  wire[46:0] T9507;
  wire[46:0] T9508;
  wire[46:0] T9509;
  wire[46:0] twiddle4_3_344_real;
  wire[46:0] T9510;
  wire[41:0] T9511;
  wire[41:0] T9512;
  wire[4:0] T9513;
  wire T9514;
  wire[46:0] T9515;
  wire[46:0] T9516;
  wire[46:0] twiddle4_3_345_real;
  wire[46:0] T9517;
  wire[42:0] T9518;
  wire[42:0] T9519;
  wire[3:0] T9520;
  wire T9521;
  wire[46:0] T9522;
  wire[46:0] T9523;
  wire T9524;
  wire[46:0] T9525;
  wire[46:0] twiddle4_3_346_real;
  wire[46:0] T9526;
  wire[42:0] T9527;
  wire[42:0] T9528;
  wire[3:0] T9529;
  wire T9530;
  wire[46:0] T9531;
  wire[46:0] T9532;
  wire[46:0] twiddle4_3_347_real;
  wire[46:0] T9533;
  wire[42:0] T9534;
  wire[42:0] T9535;
  wire[3:0] T9536;
  wire T9537;
  wire[46:0] T9538;
  wire[46:0] T9539;
  wire T9540;
  wire T9541;
  wire[46:0] T9542;
  wire[46:0] T9543;
  wire[46:0] twiddle4_3_348_real;
  wire[46:0] T9544;
  wire[42:0] T9545;
  wire[42:0] T9546;
  wire[3:0] T9547;
  wire T9548;
  wire[46:0] T9549;
  wire[46:0] T9550;
  wire[46:0] twiddle4_3_349_real;
  wire[46:0] T9551;
  wire[43:0] T9552;
  wire[43:0] T9553;
  wire[2:0] T9554;
  wire T9555;
  wire[46:0] T9556;
  wire[46:0] T9557;
  wire T9558;
  wire[46:0] T9559;
  wire[46:0] twiddle4_3_350_real;
  wire[46:0] T9560;
  wire[43:0] T9561;
  wire[43:0] T9562;
  wire[2:0] T9563;
  wire T9564;
  wire[46:0] T9565;
  wire[46:0] T9566;
  wire[46:0] twiddle4_3_351_real;
  wire[46:0] T9567;
  wire[43:0] T9568;
  wire[43:0] T9569;
  wire[2:0] T9570;
  wire T9571;
  wire[46:0] T9572;
  wire[46:0] T9573;
  wire T9574;
  wire T9575;
  wire T9576;
  wire T9577;
  wire T9578;
  wire[46:0] T9579;
  wire[46:0] T9580;
  wire[46:0] T9581;
  wire[46:0] T9582;
  wire[46:0] T9583;
  wire[46:0] twiddle4_3_352_real;
  wire[46:0] T9584;
  wire[43:0] T9585;
  wire[43:0] T9586;
  wire[2:0] T9587;
  wire T9588;
  wire[46:0] T9589;
  wire[46:0] T9590;
  wire[46:0] twiddle4_3_353_real;
  wire[46:0] T9591;
  wire[43:0] T9592;
  wire[43:0] T9593;
  wire[2:0] T9594;
  wire T9595;
  wire[46:0] T9596;
  wire[46:0] T9597;
  wire T9598;
  wire[46:0] T9599;
  wire[46:0] twiddle4_3_354_real;
  wire[46:0] T9600;
  wire[43:0] T9601;
  wire[43:0] T9602;
  wire[2:0] T9603;
  wire T9604;
  wire[46:0] T9605;
  wire[46:0] T9606;
  wire[46:0] twiddle4_3_355_real;
  wire[46:0] T9607;
  wire[44:0] T9608;
  wire[44:0] T9609;
  wire[1:0] T9610;
  wire T9611;
  wire[46:0] T9612;
  wire[46:0] T9613;
  wire T9614;
  wire T9615;
  wire[46:0] T9616;
  wire[46:0] T9617;
  wire[46:0] twiddle4_3_356_real;
  wire[46:0] T9618;
  wire[44:0] T9619;
  wire[44:0] T9620;
  wire[1:0] T9621;
  wire T9622;
  wire[46:0] T9623;
  wire[46:0] T9624;
  wire[46:0] twiddle4_3_357_real;
  wire[46:0] T9625;
  wire[44:0] T9626;
  wire[44:0] T9627;
  wire[1:0] T9628;
  wire T9629;
  wire[46:0] T9630;
  wire[46:0] T9631;
  wire T9632;
  wire[46:0] T9633;
  wire[46:0] twiddle4_3_358_real;
  wire[46:0] T9634;
  wire[44:0] T9635;
  wire[44:0] T9636;
  wire[1:0] T9637;
  wire T9638;
  wire[46:0] T9639;
  wire[46:0] T9640;
  wire[46:0] twiddle4_3_359_real;
  wire[46:0] T9641;
  wire[44:0] T9642;
  wire[44:0] T9643;
  wire[1:0] T9644;
  wire T9645;
  wire[46:0] T9646;
  wire[46:0] T9647;
  wire T9648;
  wire T9649;
  wire T9650;
  wire[46:0] T9651;
  wire[46:0] T9652;
  wire[46:0] T9653;
  wire[46:0] twiddle4_3_360_real;
  wire[46:0] T9654;
  wire[44:0] T9655;
  wire[44:0] T9656;
  wire[1:0] T9657;
  wire T9658;
  wire[46:0] T9659;
  wire[46:0] T9660;
  wire[46:0] twiddle4_3_361_real;
  wire[46:0] T9661;
  wire[44:0] T9662;
  wire[44:0] T9663;
  wire[1:0] T9664;
  wire T9665;
  wire[46:0] T9666;
  wire[46:0] T9667;
  wire T9668;
  wire[46:0] T9669;
  wire[46:0] twiddle4_3_362_real;
  wire[46:0] T9670;
  wire[44:0] T9671;
  wire[44:0] T9672;
  wire[1:0] T9673;
  wire T9674;
  wire[46:0] T9675;
  wire[46:0] T9676;
  wire[46:0] twiddle4_3_363_real;
  wire[46:0] T9677;
  wire[44:0] T9678;
  wire[44:0] T9679;
  wire[1:0] T9680;
  wire T9681;
  wire[46:0] T9682;
  wire[46:0] T9683;
  wire T9684;
  wire T9685;
  wire[46:0] T9686;
  wire[46:0] T9687;
  wire[46:0] twiddle4_3_364_real;
  wire[46:0] T9688;
  wire[44:0] T9689;
  wire[44:0] T9690;
  wire[1:0] T9691;
  wire T9692;
  wire[46:0] T9693;
  wire[46:0] T9694;
  wire[46:0] twiddle4_3_365_real;
  wire[46:0] T9695;
  wire[44:0] T9696;
  wire[44:0] T9697;
  wire[1:0] T9698;
  wire T9699;
  wire[46:0] T9700;
  wire[46:0] T9701;
  wire T9702;
  wire[46:0] T9703;
  wire[46:0] twiddle4_3_366_real;
  wire[46:0] T9704;
  wire[44:0] T9705;
  wire[44:0] T9706;
  wire[1:0] T9707;
  wire T9708;
  wire[46:0] T9709;
  wire[46:0] T9710;
  wire[46:0] twiddle4_3_367_real;
  wire[46:0] T9711;
  wire[44:0] T9712;
  wire[44:0] T9713;
  wire[1:0] T9714;
  wire T9715;
  wire[46:0] T9716;
  wire[46:0] T9717;
  wire T9718;
  wire T9719;
  wire T9720;
  wire T9721;
  wire[46:0] T9722;
  wire[46:0] T9723;
  wire[46:0] T9724;
  wire[46:0] T9725;
  wire[46:0] twiddle4_3_368_real;
  wire[46:0] T9726;
  wire[44:0] T9727;
  wire[44:0] T9728;
  wire[1:0] T9729;
  wire T9730;
  wire[46:0] T9731;
  wire[46:0] T9732;
  wire[46:0] twiddle4_3_369_real;
  wire[46:0] T9733;
  wire[45:0] T9734;
  wire[45:0] T9735;
  wire T9736;
  wire[46:0] T9737;
  wire[46:0] T9738;
  wire T9739;
  wire[46:0] T9740;
  wire[46:0] twiddle4_3_370_real;
  wire[46:0] T9741;
  wire[45:0] T9742;
  wire[45:0] T9743;
  wire T9744;
  wire[46:0] T9745;
  wire[46:0] T9746;
  wire[46:0] twiddle4_3_371_real;
  wire[46:0] T9747;
  wire[45:0] T9748;
  wire[45:0] T9749;
  wire T9750;
  wire[46:0] T9751;
  wire[46:0] T9752;
  wire T9753;
  wire T9754;
  wire[46:0] T9755;
  wire[46:0] T9756;
  wire[46:0] twiddle4_3_372_real;
  wire[46:0] T9757;
  wire[45:0] T9758;
  wire[45:0] T9759;
  wire T9760;
  wire[46:0] T9761;
  wire[46:0] T9762;
  wire[46:0] twiddle4_3_373_real;
  wire[46:0] T9763;
  wire[45:0] T9764;
  wire[45:0] T9765;
  wire T9766;
  wire[46:0] T9767;
  wire[46:0] T9768;
  wire T9769;
  wire[46:0] T9770;
  wire[46:0] twiddle4_3_374_real;
  wire[46:0] T9771;
  wire[45:0] T9772;
  wire[45:0] T9773;
  wire T9774;
  wire[46:0] T9775;
  wire[46:0] T9776;
  wire[46:0] twiddle4_3_375_real;
  wire[46:0] T9777;
  wire[45:0] T9778;
  wire[45:0] T9779;
  wire T9780;
  wire[46:0] T9781;
  wire[46:0] T9782;
  wire T9783;
  wire T9784;
  wire T9785;
  wire[46:0] T9786;
  wire[46:0] T9787;
  wire[46:0] T9788;
  wire[46:0] twiddle4_3_376_real;
  wire[46:0] T9789;
  wire[45:0] T9790;
  wire[45:0] T9791;
  wire T9792;
  wire[46:0] T9793;
  wire[46:0] T9794;
  wire[46:0] twiddle4_3_377_real;
  wire[46:0] T9795;
  wire[45:0] T9796;
  wire[45:0] T9797;
  wire T9798;
  wire[46:0] T9799;
  wire[46:0] T9800;
  wire T9801;
  wire[46:0] T9802;
  wire[46:0] twiddle4_3_378_real;
  wire[46:0] T9803;
  wire[45:0] T9804;
  wire[45:0] T9805;
  wire T9806;
  wire[46:0] T9807;
  wire[46:0] T9808;
  wire[46:0] twiddle4_3_379_real;
  wire[46:0] T9809;
  wire[45:0] T9810;
  wire[45:0] T9811;
  wire T9812;
  wire[46:0] T9813;
  wire[46:0] T9814;
  wire T9815;
  wire T9816;
  wire[46:0] T9817;
  wire[46:0] T9818;
  wire[46:0] twiddle4_3_380_real;
  wire[46:0] T9819;
  wire[45:0] T9820;
  wire[45:0] T9821;
  wire T9822;
  wire[46:0] T9823;
  wire[46:0] T9824;
  wire[46:0] twiddle4_3_381_real;
  wire[46:0] T9825;
  wire[45:0] T9826;
  wire[45:0] T9827;
  wire T9828;
  wire[46:0] T9829;
  wire[46:0] T9830;
  wire T9831;
  wire[46:0] T9832;
  wire[46:0] twiddle4_3_382_real;
  wire[46:0] T9833;
  wire[45:0] T9834;
  wire[45:0] T9835;
  wire T9836;
  wire[46:0] T9837;
  wire[46:0] T9838;
  wire[46:0] twiddle4_3_383_real;
  wire[46:0] T9839;
  wire[45:0] T9840;
  wire[45:0] T9841;
  wire T9842;
  wire[46:0] T9843;
  wire[46:0] T9844;
  wire T9845;
  wire T9846;
  wire T9847;
  wire T9848;
  wire T9849;
  wire T9850;
  wire T9851;
  wire[46:0] T9852;
  wire[46:0] T9853;
  wire[46:0] T9854;
  wire[46:0] T9855;
  wire[46:0] T9856;
  wire[46:0] T9857;
  wire[46:0] T9858;
  wire[46:0] twiddle4_3_384_real;
  wire[46:0] T9859;
  wire[45:0] T9860;
  wire[45:0] T9861;
  wire T9862;
  wire[46:0] T9863;
  wire[46:0] T9864;
  wire[46:0] twiddle4_3_385_real;
  wire[46:0] T9865;
  wire[45:0] T9866;
  wire[45:0] T9867;
  wire T9868;
  wire[46:0] T9869;
  wire[46:0] T9870;
  wire T9871;
  wire[46:0] T9872;
  wire[46:0] twiddle4_3_386_real;
  wire[46:0] T9873;
  wire[45:0] T9874;
  wire[45:0] T9875;
  wire T9876;
  wire[46:0] T9877;
  wire[46:0] T9878;
  wire[46:0] twiddle4_3_387_real;
  wire[46:0] T9879;
  wire[45:0] T9880;
  wire[45:0] T9881;
  wire T9882;
  wire[46:0] T9883;
  wire[46:0] T9884;
  wire T9885;
  wire T9886;
  wire[46:0] T9887;
  wire[46:0] T9888;
  wire[46:0] twiddle4_3_388_real;
  wire[46:0] T9889;
  wire[45:0] T9890;
  wire[45:0] T9891;
  wire T9892;
  wire[46:0] T9893;
  wire[46:0] T9894;
  wire[46:0] twiddle4_3_389_real;
  wire[46:0] T9895;
  wire[45:0] T9896;
  wire[45:0] T9897;
  wire T9898;
  wire[46:0] T9899;
  wire[46:0] T9900;
  wire T9901;
  wire[46:0] T9902;
  wire[46:0] twiddle4_3_390_real;
  wire[46:0] T9903;
  wire[45:0] T9904;
  wire[45:0] T9905;
  wire T9906;
  wire[46:0] T9907;
  wire[46:0] T9908;
  wire[46:0] twiddle4_3_391_real;
  wire[46:0] T9909;
  wire[45:0] T9910;
  wire[45:0] T9911;
  wire T9912;
  wire[46:0] T9913;
  wire[46:0] T9914;
  wire T9915;
  wire T9916;
  wire T9917;
  wire[46:0] T9918;
  wire[46:0] T9919;
  wire[46:0] T9920;
  wire[46:0] twiddle4_3_392_real;
  wire[46:0] T9921;
  wire[45:0] T9922;
  wire[45:0] T9923;
  wire T9924;
  wire[46:0] T9925;
  wire[46:0] T9926;
  wire[46:0] twiddle4_3_393_real;
  wire[46:0] T9927;
  wire[45:0] T9928;
  wire[45:0] T9929;
  wire T9930;
  wire[46:0] T9931;
  wire[46:0] T9932;
  wire T9933;
  wire[46:0] T9934;
  wire[46:0] twiddle4_3_394_real;
  wire[46:0] T9935;
  wire[45:0] T9936;
  wire[45:0] T9937;
  wire T9938;
  wire[46:0] T9939;
  wire[46:0] T9940;
  wire[46:0] twiddle4_3_395_real;
  wire[46:0] T9941;
  wire[45:0] T9942;
  wire[45:0] T9943;
  wire T9944;
  wire[46:0] T9945;
  wire[46:0] T9946;
  wire T9947;
  wire T9948;
  wire[46:0] T9949;
  wire[46:0] T9950;
  wire[46:0] twiddle4_3_396_real;
  wire[46:0] T9951;
  wire[45:0] T9952;
  wire[45:0] T9953;
  wire T9954;
  wire[46:0] T9955;
  wire[46:0] T9956;
  wire[46:0] twiddle4_3_397_real;
  wire[46:0] T9957;
  wire[45:0] T9958;
  wire[45:0] T9959;
  wire T9960;
  wire[46:0] T9961;
  wire[46:0] T9962;
  wire T9963;
  wire[46:0] T9964;
  wire[46:0] twiddle4_3_398_real;
  wire[46:0] T9965;
  wire[45:0] T9966;
  wire[45:0] T9967;
  wire T9968;
  wire[46:0] T9969;
  wire[46:0] T9970;
  wire[46:0] twiddle4_3_399_real;
  wire[46:0] T9971;
  wire[46:0] T9972;
  wire[46:0] T9973;
  wire[46:0] T9974;
  wire T9975;
  wire T9976;
  wire T9977;
  wire T9978;
  wire[46:0] T9979;
  wire[46:0] T9980;
  wire[46:0] T9981;
  wire[46:0] T9982;
  wire[46:0] twiddle4_3_400_real;
  wire[46:0] T9983;
  wire[46:0] T9984;
  wire[46:0] T9985;
  wire[46:0] T9986;
  wire[46:0] twiddle4_3_401_real;
  wire[46:0] T9987;
  wire[46:0] T9988;
  wire[46:0] T9989;
  wire[46:0] T9990;
  wire T9991;
  wire[46:0] T9992;
  wire[46:0] twiddle4_3_402_real;
  wire[46:0] T9993;
  wire[46:0] T9994;
  wire[46:0] T9995;
  wire[46:0] T9996;
  wire[46:0] twiddle4_3_403_real;
  wire[46:0] T9997;
  wire[46:0] T9998;
  wire[46:0] T9999;
  wire[46:0] T10000;
  wire T10001;
  wire T10002;
  wire[46:0] T10003;
  wire[46:0] T10004;
  wire[46:0] twiddle4_3_404_real;
  wire[46:0] T10005;
  wire[46:0] T10006;
  wire[46:0] T10007;
  wire[46:0] T10008;
  wire[46:0] twiddle4_3_405_real;
  wire[46:0] T10009;
  wire[46:0] T10010;
  wire[46:0] T10011;
  wire[46:0] T10012;
  wire T10013;
  wire[46:0] T10014;
  wire[46:0] twiddle4_3_406_real;
  wire[46:0] T10015;
  wire[46:0] T10016;
  wire[46:0] T10017;
  wire[46:0] T10018;
  wire[46:0] twiddle4_3_407_real;
  wire[46:0] T10019;
  wire[46:0] T10020;
  wire[46:0] T10021;
  wire[46:0] T10022;
  wire T10023;
  wire T10024;
  wire T10025;
  wire[46:0] T10026;
  wire[46:0] T10027;
  wire[46:0] T10028;
  wire[46:0] twiddle4_3_408_real;
  wire[46:0] T10029;
  wire[46:0] T10030;
  wire[46:0] T10031;
  wire[46:0] T10032;
  wire[46:0] twiddle4_3_409_real;
  wire[46:0] T10033;
  wire[46:0] T10034;
  wire[46:0] T10035;
  wire[46:0] T10036;
  wire T10037;
  wire[46:0] T10038;
  wire[46:0] twiddle4_3_410_real;
  wire[46:0] T10039;
  wire[46:0] T10040;
  wire[46:0] T10041;
  wire[46:0] T10042;
  wire[46:0] twiddle4_3_411_real;
  wire[46:0] T10043;
  wire[46:0] T10044;
  wire[46:0] T10045;
  wire[46:0] T10046;
  wire T10047;
  wire T10048;
  wire[46:0] T10049;
  wire[46:0] T10050;
  wire[46:0] twiddle4_3_412_real;
  wire[46:0] T10051;
  wire[46:0] T10052;
  wire[46:0] T10053;
  wire[46:0] T10054;
  wire[46:0] twiddle4_3_413_real;
  wire[46:0] T10055;
  wire[46:0] T10056;
  wire[46:0] T10057;
  wire[46:0] T10058;
  wire T10059;
  wire[46:0] T10060;
  wire[46:0] twiddle4_3_414_real;
  wire[46:0] T10061;
  wire[46:0] T10062;
  wire[46:0] T10063;
  wire[46:0] T10064;
  wire[46:0] twiddle4_3_415_real;
  wire[46:0] T10065;
  wire[46:0] T10066;
  wire[46:0] T10067;
  wire[46:0] T10068;
  wire T10069;
  wire T10070;
  wire T10071;
  wire T10072;
  wire T10073;
  wire[46:0] T10074;
  wire[46:0] T10075;
  wire[46:0] T10076;
  wire[46:0] T10077;
  wire[46:0] T10078;
  wire[46:0] twiddle4_3_416_real;
  wire[46:0] T10079;
  wire[46:0] T10080;
  wire[46:0] T10081;
  wire[46:0] T10082;
  wire[46:0] twiddle4_3_417_real;
  wire[46:0] T10083;
  wire[46:0] T10084;
  wire[46:0] T10085;
  wire[46:0] T10086;
  wire T10087;
  wire[46:0] T10088;
  wire[46:0] twiddle4_3_418_real;
  wire[46:0] T10089;
  wire[46:0] T10090;
  wire[46:0] T10091;
  wire[46:0] T10092;
  wire[46:0] twiddle4_3_419_real;
  wire[46:0] T10093;
  wire[46:0] T10094;
  wire[46:0] T10095;
  wire[46:0] T10096;
  wire T10097;
  wire T10098;
  wire[46:0] T10099;
  wire[46:0] T10100;
  wire[46:0] twiddle4_3_420_real;
  wire[46:0] T10101;
  wire[46:0] T10102;
  wire[46:0] T10103;
  wire[46:0] T10104;
  wire[46:0] twiddle4_3_421_real;
  wire[46:0] T10105;
  wire[46:0] T10106;
  wire[46:0] T10107;
  wire[46:0] T10108;
  wire T10109;
  wire[46:0] T10110;
  wire[46:0] twiddle4_3_422_real;
  wire[46:0] T10111;
  wire[46:0] T10112;
  wire[46:0] T10113;
  wire[46:0] T10114;
  wire[46:0] twiddle4_3_423_real;
  wire[46:0] T10115;
  wire[46:0] T10116;
  wire[46:0] T10117;
  wire[46:0] T10118;
  wire T10119;
  wire T10120;
  wire T10121;
  wire[46:0] T10122;
  wire[46:0] T10123;
  wire[46:0] T10124;
  wire[46:0] twiddle4_3_424_real;
  wire[46:0] T10125;
  wire[46:0] T10126;
  wire[46:0] T10127;
  wire[46:0] T10128;
  wire[46:0] twiddle4_3_425_real;
  wire[46:0] T10129;
  wire[46:0] T10130;
  wire[46:0] T10131;
  wire[46:0] T10132;
  wire T10133;
  wire[46:0] T10134;
  wire[46:0] twiddle4_3_426_real;
  wire[46:0] T10135;
  wire[46:0] T10136;
  wire[46:0] T10137;
  wire[46:0] T10138;
  wire[46:0] twiddle4_3_427_real;
  wire[46:0] T10139;
  wire[46:0] T10140;
  wire[46:0] T10141;
  wire[46:0] T10142;
  wire T10143;
  wire T10144;
  wire[46:0] T10145;
  wire[46:0] T10146;
  wire[46:0] twiddle4_3_428_real;
  wire[46:0] T10147;
  wire[46:0] T10148;
  wire[46:0] T10149;
  wire[46:0] T10150;
  wire[46:0] twiddle4_3_429_real;
  wire[46:0] T10151;
  wire[46:0] T10152;
  wire[46:0] T10153;
  wire[46:0] T10154;
  wire T10155;
  wire[46:0] T10156;
  wire[46:0] twiddle4_3_430_real;
  wire[46:0] T10157;
  wire[46:0] T10158;
  wire[46:0] T10159;
  wire[46:0] T10160;
  wire[46:0] twiddle4_3_431_real;
  wire[46:0] T10161;
  wire[46:0] T10162;
  wire[46:0] T10163;
  wire[46:0] T10164;
  wire T10165;
  wire T10166;
  wire T10167;
  wire T10168;
  wire[46:0] T10169;
  wire[46:0] T10170;
  wire[46:0] T10171;
  wire[46:0] T10172;
  wire[46:0] twiddle4_3_432_real;
  wire[46:0] T10173;
  wire[46:0] T10174;
  wire[46:0] T10175;
  wire[46:0] T10176;
  wire[46:0] twiddle4_3_433_real;
  wire[46:0] T10177;
  wire[46:0] T10178;
  wire[46:0] T10179;
  wire[46:0] T10180;
  wire T10181;
  wire[46:0] T10182;
  wire[46:0] twiddle4_3_434_real;
  wire[46:0] T10183;
  wire[46:0] T10184;
  wire[46:0] T10185;
  wire[46:0] T10186;
  wire[46:0] twiddle4_3_435_real;
  wire[46:0] T10187;
  wire[46:0] T10188;
  wire[46:0] T10189;
  wire[46:0] T10190;
  wire T10191;
  wire T10192;
  wire[46:0] T10193;
  wire[46:0] T10194;
  wire[46:0] twiddle4_3_436_real;
  wire[46:0] T10195;
  wire[46:0] T10196;
  wire[46:0] T10197;
  wire[46:0] T10198;
  wire[46:0] twiddle4_3_437_real;
  wire[46:0] T10199;
  wire[46:0] T10200;
  wire[46:0] T10201;
  wire[46:0] T10202;
  wire T10203;
  wire[46:0] T10204;
  wire[46:0] twiddle4_3_438_real;
  wire[46:0] T10205;
  wire[46:0] T10206;
  wire[46:0] T10207;
  wire[46:0] T10208;
  wire[46:0] twiddle4_3_439_real;
  wire[46:0] T10209;
  wire[46:0] T10210;
  wire[46:0] T10211;
  wire[46:0] T10212;
  wire T10213;
  wire T10214;
  wire T10215;
  wire[46:0] T10216;
  wire[46:0] T10217;
  wire[46:0] T10218;
  wire[46:0] twiddle4_3_440_real;
  wire[46:0] T10219;
  wire[46:0] T10220;
  wire[46:0] T10221;
  wire[46:0] T10222;
  wire[46:0] twiddle4_3_441_real;
  wire[46:0] T10223;
  wire[46:0] T10224;
  wire[46:0] T10225;
  wire[46:0] T10226;
  wire T10227;
  wire[46:0] T10228;
  wire[46:0] twiddle4_3_442_real;
  wire[46:0] T10229;
  wire[46:0] T10230;
  wire[46:0] T10231;
  wire[46:0] T10232;
  wire[46:0] twiddle4_3_443_real;
  wire[46:0] T10233;
  wire[46:0] T10234;
  wire[46:0] T10235;
  wire[46:0] T10236;
  wire T10237;
  wire T10238;
  wire[46:0] T10239;
  wire[46:0] T10240;
  wire[46:0] twiddle4_3_444_real;
  wire[46:0] T10241;
  wire[46:0] T10242;
  wire[46:0] T10243;
  wire[46:0] T10244;
  wire[46:0] twiddle4_3_445_real;
  wire[46:0] T10245;
  wire[46:0] T10246;
  wire[46:0] T10247;
  wire[46:0] T10248;
  wire T10249;
  wire[46:0] T10250;
  wire[46:0] twiddle4_3_446_real;
  wire[46:0] T10251;
  wire[46:0] T10252;
  wire[46:0] T10253;
  wire[46:0] T10254;
  wire[46:0] twiddle4_3_447_real;
  wire[46:0] T10255;
  wire[46:0] T10256;
  wire[46:0] T10257;
  wire[46:0] T10258;
  wire T10259;
  wire T10260;
  wire T10261;
  wire T10262;
  wire T10263;
  wire T10264;
  wire[46:0] T10265;
  wire[46:0] T10266;
  wire[46:0] T10267;
  wire[46:0] T10268;
  wire[46:0] T10269;
  wire[46:0] T10270;
  wire[46:0] twiddle4_3_448_real;
  wire[46:0] T10271;
  wire[46:0] T10272;
  wire[46:0] T10273;
  wire[46:0] T10274;
  wire[46:0] twiddle4_3_449_real;
  wire[46:0] T10275;
  wire[46:0] T10276;
  wire[46:0] T10277;
  wire[46:0] T10278;
  wire T10279;
  wire[46:0] T10280;
  wire[46:0] twiddle4_3_450_real;
  wire[46:0] T10281;
  wire[46:0] T10282;
  wire[46:0] T10283;
  wire[46:0] T10284;
  wire[46:0] twiddle4_3_451_real;
  wire[46:0] T10285;
  wire[46:0] T10286;
  wire[46:0] T10287;
  wire[46:0] T10288;
  wire T10289;
  wire T10290;
  wire[46:0] T10291;
  wire[46:0] T10292;
  wire[46:0] twiddle4_3_452_real;
  wire[46:0] T10293;
  wire[46:0] T10294;
  wire[46:0] T10295;
  wire[46:0] T10296;
  wire[46:0] twiddle4_3_453_real;
  wire[46:0] T10297;
  wire[46:0] T10298;
  wire[46:0] T10299;
  wire[46:0] T10300;
  wire T10301;
  wire[46:0] T10302;
  wire[46:0] twiddle4_3_454_real;
  wire[46:0] T10303;
  wire[46:0] T10304;
  wire[46:0] T10305;
  wire[46:0] T10306;
  wire[46:0] twiddle4_3_455_real;
  wire[46:0] T10307;
  wire[46:0] T10308;
  wire[46:0] T10309;
  wire[46:0] T10310;
  wire T10311;
  wire T10312;
  wire T10313;
  wire[46:0] T10314;
  wire[46:0] T10315;
  wire[46:0] T10316;
  wire[46:0] twiddle4_3_456_real;
  wire[46:0] T10317;
  wire[46:0] T10318;
  wire[46:0] T10319;
  wire[45:0] T10320;
  wire[45:0] T10321;
  wire T10322;
  wire[46:0] twiddle4_3_457_real;
  wire[46:0] T10323;
  wire[46:0] T10324;
  wire[46:0] T10325;
  wire[45:0] T10326;
  wire[45:0] T10327;
  wire T10328;
  wire T10329;
  wire[46:0] T10330;
  wire[46:0] twiddle4_3_458_real;
  wire[46:0] T10331;
  wire[46:0] T10332;
  wire[46:0] T10333;
  wire[45:0] T10334;
  wire[45:0] T10335;
  wire T10336;
  wire[46:0] twiddle4_3_459_real;
  wire[46:0] T10337;
  wire[46:0] T10338;
  wire[46:0] T10339;
  wire[45:0] T10340;
  wire[45:0] T10341;
  wire T10342;
  wire T10343;
  wire T10344;
  wire[46:0] T10345;
  wire[46:0] T10346;
  wire[46:0] twiddle4_3_460_real;
  wire[46:0] T10347;
  wire[46:0] T10348;
  wire[46:0] T10349;
  wire[45:0] T10350;
  wire[45:0] T10351;
  wire T10352;
  wire[46:0] twiddle4_3_461_real;
  wire[46:0] T10353;
  wire[46:0] T10354;
  wire[46:0] T10355;
  wire[45:0] T10356;
  wire[45:0] T10357;
  wire T10358;
  wire T10359;
  wire[46:0] T10360;
  wire[46:0] twiddle4_3_462_real;
  wire[46:0] T10361;
  wire[46:0] T10362;
  wire[46:0] T10363;
  wire[45:0] T10364;
  wire[45:0] T10365;
  wire T10366;
  wire[46:0] twiddle4_3_463_real;
  wire[46:0] T10367;
  wire[46:0] T10368;
  wire[46:0] T10369;
  wire[45:0] T10370;
  wire[45:0] T10371;
  wire T10372;
  wire T10373;
  wire T10374;
  wire T10375;
  wire T10376;
  wire[46:0] T10377;
  wire[46:0] T10378;
  wire[46:0] T10379;
  wire[46:0] T10380;
  wire[46:0] twiddle4_3_464_real;
  wire[46:0] T10381;
  wire[46:0] T10382;
  wire[46:0] T10383;
  wire[45:0] T10384;
  wire[45:0] T10385;
  wire T10386;
  wire[46:0] twiddle4_3_465_real;
  wire[46:0] T10387;
  wire[46:0] T10388;
  wire[46:0] T10389;
  wire[45:0] T10390;
  wire[45:0] T10391;
  wire T10392;
  wire T10393;
  wire[46:0] T10394;
  wire[46:0] twiddle4_3_466_real;
  wire[46:0] T10395;
  wire[46:0] T10396;
  wire[46:0] T10397;
  wire[45:0] T10398;
  wire[45:0] T10399;
  wire T10400;
  wire[46:0] twiddle4_3_467_real;
  wire[46:0] T10401;
  wire[46:0] T10402;
  wire[46:0] T10403;
  wire[45:0] T10404;
  wire[45:0] T10405;
  wire T10406;
  wire T10407;
  wire T10408;
  wire[46:0] T10409;
  wire[46:0] T10410;
  wire[46:0] twiddle4_3_468_real;
  wire[46:0] T10411;
  wire[46:0] T10412;
  wire[46:0] T10413;
  wire[45:0] T10414;
  wire[45:0] T10415;
  wire T10416;
  wire[46:0] twiddle4_3_469_real;
  wire[46:0] T10417;
  wire[46:0] T10418;
  wire[46:0] T10419;
  wire[45:0] T10420;
  wire[45:0] T10421;
  wire T10422;
  wire T10423;
  wire[46:0] T10424;
  wire[46:0] twiddle4_3_470_real;
  wire[46:0] T10425;
  wire[46:0] T10426;
  wire[46:0] T10427;
  wire[45:0] T10428;
  wire[45:0] T10429;
  wire T10430;
  wire[46:0] twiddle4_3_471_real;
  wire[46:0] T10431;
  wire[46:0] T10432;
  wire[46:0] T10433;
  wire[45:0] T10434;
  wire[45:0] T10435;
  wire T10436;
  wire T10437;
  wire T10438;
  wire T10439;
  wire[46:0] T10440;
  wire[46:0] T10441;
  wire[46:0] T10442;
  wire[46:0] twiddle4_3_472_real;
  wire[46:0] T10443;
  wire[46:0] T10444;
  wire[46:0] T10445;
  wire[45:0] T10446;
  wire[45:0] T10447;
  wire T10448;
  wire[46:0] twiddle4_3_473_real;
  wire[46:0] T10449;
  wire[46:0] T10450;
  wire[46:0] T10451;
  wire[45:0] T10452;
  wire[45:0] T10453;
  wire T10454;
  wire T10455;
  wire[46:0] T10456;
  wire[46:0] twiddle4_3_474_real;
  wire[46:0] T10457;
  wire[46:0] T10458;
  wire[46:0] T10459;
  wire[45:0] T10460;
  wire[45:0] T10461;
  wire T10462;
  wire[46:0] twiddle4_3_475_real;
  wire[46:0] T10463;
  wire[46:0] T10464;
  wire[46:0] T10465;
  wire[45:0] T10466;
  wire[45:0] T10467;
  wire T10468;
  wire T10469;
  wire T10470;
  wire[46:0] T10471;
  wire[46:0] T10472;
  wire[46:0] twiddle4_3_476_real;
  wire[46:0] T10473;
  wire[46:0] T10474;
  wire[46:0] T10475;
  wire[45:0] T10476;
  wire[45:0] T10477;
  wire T10478;
  wire[46:0] twiddle4_3_477_real;
  wire[46:0] T10479;
  wire[46:0] T10480;
  wire[46:0] T10481;
  wire[45:0] T10482;
  wire[45:0] T10483;
  wire T10484;
  wire T10485;
  wire[46:0] T10486;
  wire[46:0] twiddle4_3_478_real;
  wire[46:0] T10487;
  wire[46:0] T10488;
  wire[46:0] T10489;
  wire[45:0] T10490;
  wire[45:0] T10491;
  wire T10492;
  wire[46:0] twiddle4_3_479_real;
  wire[46:0] T10493;
  wire[46:0] T10494;
  wire[46:0] T10495;
  wire[45:0] T10496;
  wire[45:0] T10497;
  wire T10498;
  wire T10499;
  wire T10500;
  wire T10501;
  wire T10502;
  wire T10503;
  wire[46:0] T10504;
  wire[46:0] T10505;
  wire[46:0] T10506;
  wire[46:0] T10507;
  wire[46:0] T10508;
  wire[46:0] twiddle4_3_480_real;
  wire[46:0] T10509;
  wire[46:0] T10510;
  wire[46:0] T10511;
  wire[45:0] T10512;
  wire[45:0] T10513;
  wire T10514;
  wire[46:0] twiddle4_3_481_real;
  wire[46:0] T10515;
  wire[46:0] T10516;
  wire[46:0] T10517;
  wire[45:0] T10518;
  wire[45:0] T10519;
  wire T10520;
  wire T10521;
  wire[46:0] T10522;
  wire[46:0] twiddle4_3_482_real;
  wire[46:0] T10523;
  wire[46:0] T10524;
  wire[46:0] T10525;
  wire[45:0] T10526;
  wire[45:0] T10527;
  wire T10528;
  wire[46:0] twiddle4_3_483_real;
  wire[46:0] T10529;
  wire[46:0] T10530;
  wire[46:0] T10531;
  wire[45:0] T10532;
  wire[45:0] T10533;
  wire T10534;
  wire T10535;
  wire T10536;
  wire[46:0] T10537;
  wire[46:0] T10538;
  wire[46:0] twiddle4_3_484_real;
  wire[46:0] T10539;
  wire[46:0] T10540;
  wire[46:0] T10541;
  wire[45:0] T10542;
  wire[45:0] T10543;
  wire T10544;
  wire[46:0] twiddle4_3_485_real;
  wire[46:0] T10545;
  wire[46:0] T10546;
  wire[46:0] T10547;
  wire[44:0] T10548;
  wire[44:0] T10549;
  wire[1:0] T10550;
  wire T10551;
  wire T10552;
  wire[46:0] T10553;
  wire[46:0] twiddle4_3_486_real;
  wire[46:0] T10554;
  wire[46:0] T10555;
  wire[46:0] T10556;
  wire[44:0] T10557;
  wire[44:0] T10558;
  wire[1:0] T10559;
  wire T10560;
  wire[46:0] twiddle4_3_487_real;
  wire[46:0] T10561;
  wire[46:0] T10562;
  wire[46:0] T10563;
  wire[44:0] T10564;
  wire[44:0] T10565;
  wire[1:0] T10566;
  wire T10567;
  wire T10568;
  wire T10569;
  wire T10570;
  wire[46:0] T10571;
  wire[46:0] T10572;
  wire[46:0] T10573;
  wire[46:0] twiddle4_3_488_real;
  wire[46:0] T10574;
  wire[46:0] T10575;
  wire[46:0] T10576;
  wire[44:0] T10577;
  wire[44:0] T10578;
  wire[1:0] T10579;
  wire T10580;
  wire[46:0] twiddle4_3_489_real;
  wire[46:0] T10581;
  wire[46:0] T10582;
  wire[46:0] T10583;
  wire[44:0] T10584;
  wire[44:0] T10585;
  wire[1:0] T10586;
  wire T10587;
  wire T10588;
  wire[46:0] T10589;
  wire[46:0] twiddle4_3_490_real;
  wire[46:0] T10590;
  wire[46:0] T10591;
  wire[46:0] T10592;
  wire[44:0] T10593;
  wire[44:0] T10594;
  wire[1:0] T10595;
  wire T10596;
  wire[46:0] twiddle4_3_491_real;
  wire[46:0] T10597;
  wire[46:0] T10598;
  wire[46:0] T10599;
  wire[44:0] T10600;
  wire[44:0] T10601;
  wire[1:0] T10602;
  wire T10603;
  wire T10604;
  wire T10605;
  wire[46:0] T10606;
  wire[46:0] T10607;
  wire[46:0] twiddle4_3_492_real;
  wire[46:0] T10608;
  wire[46:0] T10609;
  wire[46:0] T10610;
  wire[44:0] T10611;
  wire[44:0] T10612;
  wire[1:0] T10613;
  wire T10614;
  wire[46:0] twiddle4_3_493_real;
  wire[46:0] T10615;
  wire[46:0] T10616;
  wire[46:0] T10617;
  wire[44:0] T10618;
  wire[44:0] T10619;
  wire[1:0] T10620;
  wire T10621;
  wire T10622;
  wire[46:0] T10623;
  wire[46:0] twiddle4_3_494_real;
  wire[46:0] T10624;
  wire[46:0] T10625;
  wire[46:0] T10626;
  wire[44:0] T10627;
  wire[44:0] T10628;
  wire[1:0] T10629;
  wire T10630;
  wire[46:0] twiddle4_3_495_real;
  wire[46:0] T10631;
  wire[46:0] T10632;
  wire[46:0] T10633;
  wire[44:0] T10634;
  wire[44:0] T10635;
  wire[1:0] T10636;
  wire T10637;
  wire T10638;
  wire T10639;
  wire T10640;
  wire T10641;
  wire[46:0] T10642;
  wire[46:0] T10643;
  wire[46:0] T10644;
  wire[46:0] T10645;
  wire[46:0] twiddle4_3_496_real;
  wire[46:0] T10646;
  wire[46:0] T10647;
  wire[46:0] T10648;
  wire[44:0] T10649;
  wire[44:0] T10650;
  wire[1:0] T10651;
  wire T10652;
  wire[46:0] twiddle4_3_497_real;
  wire[46:0] T10653;
  wire[46:0] T10654;
  wire[46:0] T10655;
  wire[44:0] T10656;
  wire[44:0] T10657;
  wire[1:0] T10658;
  wire T10659;
  wire T10660;
  wire[46:0] T10661;
  wire[46:0] twiddle4_3_498_real;
  wire[46:0] T10662;
  wire[46:0] T10663;
  wire[46:0] T10664;
  wire[44:0] T10665;
  wire[44:0] T10666;
  wire[1:0] T10667;
  wire T10668;
  wire[46:0] twiddle4_3_499_real;
  wire[46:0] T10669;
  wire[46:0] T10670;
  wire[46:0] T10671;
  wire[43:0] T10672;
  wire[43:0] T10673;
  wire[2:0] T10674;
  wire T10675;
  wire T10676;
  wire T10677;
  wire[46:0] T10678;
  wire[46:0] T10679;
  wire[46:0] twiddle4_3_500_real;
  wire[46:0] T10680;
  wire[46:0] T10681;
  wire[46:0] T10682;
  wire[43:0] T10683;
  wire[43:0] T10684;
  wire[2:0] T10685;
  wire T10686;
  wire[46:0] twiddle4_3_501_real;
  wire[46:0] T10687;
  wire[46:0] T10688;
  wire[46:0] T10689;
  wire[43:0] T10690;
  wire[43:0] T10691;
  wire[2:0] T10692;
  wire T10693;
  wire T10694;
  wire[46:0] T10695;
  wire[46:0] twiddle4_3_502_real;
  wire[46:0] T10696;
  wire[46:0] T10697;
  wire[46:0] T10698;
  wire[43:0] T10699;
  wire[43:0] T10700;
  wire[2:0] T10701;
  wire T10702;
  wire[46:0] twiddle4_3_503_real;
  wire[46:0] T10703;
  wire[46:0] T10704;
  wire[46:0] T10705;
  wire[43:0] T10706;
  wire[43:0] T10707;
  wire[2:0] T10708;
  wire T10709;
  wire T10710;
  wire T10711;
  wire T10712;
  wire[46:0] T10713;
  wire[46:0] T10714;
  wire[46:0] T10715;
  wire[46:0] twiddle4_3_504_real;
  wire[46:0] T10716;
  wire[46:0] T10717;
  wire[46:0] T10718;
  wire[43:0] T10719;
  wire[43:0] T10720;
  wire[2:0] T10721;
  wire T10722;
  wire[46:0] twiddle4_3_505_real;
  wire[46:0] T10723;
  wire[46:0] T10724;
  wire[46:0] T10725;
  wire[43:0] T10726;
  wire[43:0] T10727;
  wire[2:0] T10728;
  wire T10729;
  wire T10730;
  wire[46:0] T10731;
  wire[46:0] twiddle4_3_506_real;
  wire[46:0] T10732;
  wire[46:0] T10733;
  wire[46:0] T10734;
  wire[42:0] T10735;
  wire[42:0] T10736;
  wire[3:0] T10737;
  wire T10738;
  wire[46:0] twiddle4_3_507_real;
  wire[46:0] T10739;
  wire[46:0] T10740;
  wire[46:0] T10741;
  wire[42:0] T10742;
  wire[42:0] T10743;
  wire[3:0] T10744;
  wire T10745;
  wire T10746;
  wire T10747;
  wire[46:0] T10748;
  wire[46:0] T10749;
  wire[46:0] twiddle4_3_508_real;
  wire[46:0] T10750;
  wire[46:0] T10751;
  wire[46:0] T10752;
  wire[42:0] T10753;
  wire[42:0] T10754;
  wire[3:0] T10755;
  wire T10756;
  wire[46:0] twiddle4_3_509_real;
  wire[46:0] T10757;
  wire[46:0] T10758;
  wire[46:0] T10759;
  wire[41:0] T10760;
  wire[41:0] T10761;
  wire[4:0] T10762;
  wire T10763;
  wire T10764;
  wire[46:0] T10765;
  wire[46:0] twiddle4_3_510_real;
  wire[46:0] T10766;
  wire[46:0] T10767;
  wire[46:0] T10768;
  wire[41:0] T10769;
  wire[41:0] T10770;
  wire[4:0] T10771;
  wire T10772;
  wire[46:0] twiddle4_3_511_real;
  wire[46:0] T10773;
  wire[46:0] T10774;
  wire[46:0] T10775;
  wire[40:0] T10776;
  wire[40:0] T10777;
  wire[5:0] T10778;
  wire T10779;
  wire T10780;
  wire T10781;
  wire T10782;
  wire T10783;
  wire T10784;
  wire T10785;
  wire T10786;
  wire T10787;
  wire T10788;
  wire T10789;
  wire[15:0] T10790;
  wire[47:0] T10791;
  wire[47:0] T10792;
  wire[47:0] T10793;
  wire[47:0] T10794;
  wire[47:0] T10795;
  wire[47:0] T10796;
  wire[47:0] T10797;
  wire[47:0] T10798;
  wire[47:0] T10799;
  wire[47:0] twiddle4_2_0_imag;
  wire[47:0] T10800;
  wire[16:0] T10801;
  wire[16:0] T10802;
  wire[30:0] T10803;
  wire T10804;
  wire[47:0] T10805;
  wire[47:0] T10806;
  wire[47:0] T10807;
  wire[46:0] twiddle4_2_1_imag;
  wire[46:0] T10808;
  wire[39:0] T10809;
  wire[39:0] T10810;
  wire[6:0] T10811;
  wire T10812;
  wire[46:0] T10813;
  wire[46:0] T10814;
  wire T10815;
  wire T10816;
  wire[8:0] T10817;
  wire[8:0] T10818;
  wire[47:0] T10819;
  wire[46:0] T10820;
  wire[46:0] twiddle4_2_2_imag;
  wire[46:0] T10821;
  wire[40:0] T10822;
  wire[40:0] T10823;
  wire[5:0] T10824;
  wire T10825;
  wire[46:0] T10826;
  wire[46:0] T10827;
  wire[46:0] twiddle4_2_3_imag;
  wire[46:0] T10828;
  wire[41:0] T10829;
  wire[41:0] T10830;
  wire[4:0] T10831;
  wire T10832;
  wire[46:0] T10833;
  wire[46:0] T10834;
  wire T10835;
  wire T10836;
  wire T10837;
  wire[47:0] T10838;
  wire[46:0] T10839;
  wire[46:0] T10840;
  wire[46:0] twiddle4_2_4_imag;
  wire[46:0] T10841;
  wire[41:0] T10842;
  wire[41:0] T10843;
  wire[4:0] T10844;
  wire T10845;
  wire[46:0] T10846;
  wire[46:0] T10847;
  wire[46:0] twiddle4_2_5_imag;
  wire[46:0] T10848;
  wire[41:0] T10849;
  wire[41:0] T10850;
  wire[4:0] T10851;
  wire T10852;
  wire[46:0] T10853;
  wire[46:0] T10854;
  wire T10855;
  wire[46:0] T10856;
  wire[46:0] twiddle4_2_6_imag;
  wire[46:0] T10857;
  wire[42:0] T10858;
  wire[42:0] T10859;
  wire[3:0] T10860;
  wire T10861;
  wire[46:0] T10862;
  wire[46:0] T10863;
  wire[46:0] twiddle4_2_7_imag;
  wire[46:0] T10864;
  wire[42:0] T10865;
  wire[42:0] T10866;
  wire[3:0] T10867;
  wire T10868;
  wire[46:0] T10869;
  wire[46:0] T10870;
  wire T10871;
  wire T10872;
  wire T10873;
  wire T10874;
  wire[47:0] T10875;
  wire[46:0] T10876;
  wire[46:0] T10877;
  wire[46:0] T10878;
  wire[46:0] twiddle4_2_8_imag;
  wire[46:0] T10879;
  wire[42:0] T10880;
  wire[42:0] T10881;
  wire[3:0] T10882;
  wire T10883;
  wire[46:0] T10884;
  wire[46:0] T10885;
  wire[46:0] twiddle4_2_9_imag;
  wire[46:0] T10886;
  wire[42:0] T10887;
  wire[42:0] T10888;
  wire[3:0] T10889;
  wire T10890;
  wire[46:0] T10891;
  wire[46:0] T10892;
  wire T10893;
  wire[46:0] T10894;
  wire[46:0] twiddle4_2_10_imag;
  wire[46:0] T10895;
  wire[42:0] T10896;
  wire[42:0] T10897;
  wire[3:0] T10898;
  wire T10899;
  wire[46:0] T10900;
  wire[46:0] T10901;
  wire[46:0] twiddle4_2_11_imag;
  wire[46:0] T10902;
  wire[43:0] T10903;
  wire[43:0] T10904;
  wire[2:0] T10905;
  wire T10906;
  wire[46:0] T10907;
  wire[46:0] T10908;
  wire T10909;
  wire T10910;
  wire[46:0] T10911;
  wire[46:0] T10912;
  wire[46:0] twiddle4_2_12_imag;
  wire[46:0] T10913;
  wire[43:0] T10914;
  wire[43:0] T10915;
  wire[2:0] T10916;
  wire T10917;
  wire[46:0] T10918;
  wire[46:0] T10919;
  wire[46:0] twiddle4_2_13_imag;
  wire[46:0] T10920;
  wire[43:0] T10921;
  wire[43:0] T10922;
  wire[2:0] T10923;
  wire T10924;
  wire[46:0] T10925;
  wire[46:0] T10926;
  wire T10927;
  wire[46:0] T10928;
  wire[46:0] twiddle4_2_14_imag;
  wire[46:0] T10929;
  wire[43:0] T10930;
  wire[43:0] T10931;
  wire[2:0] T10932;
  wire T10933;
  wire[46:0] T10934;
  wire[46:0] T10935;
  wire[46:0] twiddle4_2_15_imag;
  wire[46:0] T10936;
  wire[43:0] T10937;
  wire[43:0] T10938;
  wire[2:0] T10939;
  wire T10940;
  wire[46:0] T10941;
  wire[46:0] T10942;
  wire T10943;
  wire T10944;
  wire T10945;
  wire T10946;
  wire T10947;
  wire[47:0] T10948;
  wire[46:0] T10949;
  wire[46:0] T10950;
  wire[46:0] T10951;
  wire[46:0] T10952;
  wire[46:0] twiddle4_2_16_imag;
  wire[46:0] T10953;
  wire[43:0] T10954;
  wire[43:0] T10955;
  wire[2:0] T10956;
  wire T10957;
  wire[46:0] T10958;
  wire[46:0] T10959;
  wire[46:0] twiddle4_2_17_imag;
  wire[46:0] T10960;
  wire[43:0] T10961;
  wire[43:0] T10962;
  wire[2:0] T10963;
  wire T10964;
  wire[46:0] T10965;
  wire[46:0] T10966;
  wire T10967;
  wire[46:0] T10968;
  wire[46:0] twiddle4_2_18_imag;
  wire[46:0] T10969;
  wire[43:0] T10970;
  wire[43:0] T10971;
  wire[2:0] T10972;
  wire T10973;
  wire[46:0] T10974;
  wire[46:0] T10975;
  wire[46:0] twiddle4_2_19_imag;
  wire[46:0] T10976;
  wire[43:0] T10977;
  wire[43:0] T10978;
  wire[2:0] T10979;
  wire T10980;
  wire[46:0] T10981;
  wire[46:0] T10982;
  wire T10983;
  wire T10984;
  wire[46:0] T10985;
  wire[46:0] T10986;
  wire[46:0] twiddle4_2_20_imag;
  wire[46:0] T10987;
  wire[43:0] T10988;
  wire[43:0] T10989;
  wire[2:0] T10990;
  wire T10991;
  wire[46:0] T10992;
  wire[46:0] T10993;
  wire[46:0] twiddle4_2_21_imag;
  wire[46:0] T10994;
  wire[44:0] T10995;
  wire[44:0] T10996;
  wire[1:0] T10997;
  wire T10998;
  wire[46:0] T10999;
  wire[46:0] T11000;
  wire T11001;
  wire[46:0] T11002;
  wire[46:0] twiddle4_2_22_imag;
  wire[46:0] T11003;
  wire[44:0] T11004;
  wire[44:0] T11005;
  wire[1:0] T11006;
  wire T11007;
  wire[46:0] T11008;
  wire[46:0] T11009;
  wire[46:0] twiddle4_2_23_imag;
  wire[46:0] T11010;
  wire[44:0] T11011;
  wire[44:0] T11012;
  wire[1:0] T11013;
  wire T11014;
  wire[46:0] T11015;
  wire[46:0] T11016;
  wire T11017;
  wire T11018;
  wire T11019;
  wire[46:0] T11020;
  wire[46:0] T11021;
  wire[46:0] T11022;
  wire[46:0] twiddle4_2_24_imag;
  wire[46:0] T11023;
  wire[44:0] T11024;
  wire[44:0] T11025;
  wire[1:0] T11026;
  wire T11027;
  wire[46:0] T11028;
  wire[46:0] T11029;
  wire[46:0] twiddle4_2_25_imag;
  wire[46:0] T11030;
  wire[44:0] T11031;
  wire[44:0] T11032;
  wire[1:0] T11033;
  wire T11034;
  wire[46:0] T11035;
  wire[46:0] T11036;
  wire T11037;
  wire[46:0] T11038;
  wire[46:0] twiddle4_2_26_imag;
  wire[46:0] T11039;
  wire[44:0] T11040;
  wire[44:0] T11041;
  wire[1:0] T11042;
  wire T11043;
  wire[46:0] T11044;
  wire[46:0] T11045;
  wire[46:0] twiddle4_2_27_imag;
  wire[46:0] T11046;
  wire[44:0] T11047;
  wire[44:0] T11048;
  wire[1:0] T11049;
  wire T11050;
  wire[46:0] T11051;
  wire[46:0] T11052;
  wire T11053;
  wire T11054;
  wire[46:0] T11055;
  wire[46:0] T11056;
  wire[46:0] twiddle4_2_28_imag;
  wire[46:0] T11057;
  wire[44:0] T11058;
  wire[44:0] T11059;
  wire[1:0] T11060;
  wire T11061;
  wire[46:0] T11062;
  wire[46:0] T11063;
  wire[46:0] twiddle4_2_29_imag;
  wire[46:0] T11064;
  wire[44:0] T11065;
  wire[44:0] T11066;
  wire[1:0] T11067;
  wire T11068;
  wire[46:0] T11069;
  wire[46:0] T11070;
  wire T11071;
  wire[46:0] T11072;
  wire[46:0] twiddle4_2_30_imag;
  wire[46:0] T11073;
  wire[44:0] T11074;
  wire[44:0] T11075;
  wire[1:0] T11076;
  wire T11077;
  wire[46:0] T11078;
  wire[46:0] T11079;
  wire[46:0] twiddle4_2_31_imag;
  wire[46:0] T11080;
  wire[44:0] T11081;
  wire[44:0] T11082;
  wire[1:0] T11083;
  wire T11084;
  wire[46:0] T11085;
  wire[46:0] T11086;
  wire T11087;
  wire T11088;
  wire T11089;
  wire T11090;
  wire T11091;
  wire T11092;
  wire[47:0] T11093;
  wire[46:0] T11094;
  wire[46:0] T11095;
  wire[46:0] T11096;
  wire[46:0] T11097;
  wire[46:0] T11098;
  wire[46:0] twiddle4_2_32_imag;
  wire[46:0] T11099;
  wire[44:0] T11100;
  wire[44:0] T11101;
  wire[1:0] T11102;
  wire T11103;
  wire[46:0] T11104;
  wire[46:0] T11105;
  wire[46:0] twiddle4_2_33_imag;
  wire[46:0] T11106;
  wire[44:0] T11107;
  wire[44:0] T11108;
  wire[1:0] T11109;
  wire T11110;
  wire[46:0] T11111;
  wire[46:0] T11112;
  wire T11113;
  wire[46:0] T11114;
  wire[46:0] twiddle4_2_34_imag;
  wire[46:0] T11115;
  wire[44:0] T11116;
  wire[44:0] T11117;
  wire[1:0] T11118;
  wire T11119;
  wire[46:0] T11120;
  wire[46:0] T11121;
  wire[46:0] twiddle4_2_35_imag;
  wire[46:0] T11122;
  wire[44:0] T11123;
  wire[44:0] T11124;
  wire[1:0] T11125;
  wire T11126;
  wire[46:0] T11127;
  wire[46:0] T11128;
  wire T11129;
  wire T11130;
  wire[46:0] T11131;
  wire[46:0] T11132;
  wire[46:0] twiddle4_2_36_imag;
  wire[46:0] T11133;
  wire[44:0] T11134;
  wire[44:0] T11135;
  wire[1:0] T11136;
  wire T11137;
  wire[46:0] T11138;
  wire[46:0] T11139;
  wire[46:0] twiddle4_2_37_imag;
  wire[46:0] T11140;
  wire[44:0] T11141;
  wire[44:0] T11142;
  wire[1:0] T11143;
  wire T11144;
  wire[46:0] T11145;
  wire[46:0] T11146;
  wire T11147;
  wire[46:0] T11148;
  wire[46:0] twiddle4_2_38_imag;
  wire[46:0] T11149;
  wire[44:0] T11150;
  wire[44:0] T11151;
  wire[1:0] T11152;
  wire T11153;
  wire[46:0] T11154;
  wire[46:0] T11155;
  wire[46:0] twiddle4_2_39_imag;
  wire[46:0] T11156;
  wire[44:0] T11157;
  wire[44:0] T11158;
  wire[1:0] T11159;
  wire T11160;
  wire[46:0] T11161;
  wire[46:0] T11162;
  wire T11163;
  wire T11164;
  wire T11165;
  wire[46:0] T11166;
  wire[46:0] T11167;
  wire[46:0] T11168;
  wire[46:0] twiddle4_2_40_imag;
  wire[46:0] T11169;
  wire[44:0] T11170;
  wire[44:0] T11171;
  wire[1:0] T11172;
  wire T11173;
  wire[46:0] T11174;
  wire[46:0] T11175;
  wire[46:0] twiddle4_2_41_imag;
  wire[46:0] T11176;
  wire[44:0] T11177;
  wire[44:0] T11178;
  wire[1:0] T11179;
  wire T11180;
  wire[46:0] T11181;
  wire[46:0] T11182;
  wire T11183;
  wire[46:0] T11184;
  wire[46:0] twiddle4_2_42_imag;
  wire[46:0] T11185;
  wire[45:0] T11186;
  wire[45:0] T11187;
  wire T11188;
  wire[46:0] T11189;
  wire[46:0] T11190;
  wire[46:0] twiddle4_2_43_imag;
  wire[46:0] T11191;
  wire[45:0] T11192;
  wire[45:0] T11193;
  wire T11194;
  wire[46:0] T11195;
  wire[46:0] T11196;
  wire T11197;
  wire T11198;
  wire[46:0] T11199;
  wire[46:0] T11200;
  wire[46:0] twiddle4_2_44_imag;
  wire[46:0] T11201;
  wire[45:0] T11202;
  wire[45:0] T11203;
  wire T11204;
  wire[46:0] T11205;
  wire[46:0] T11206;
  wire[46:0] twiddle4_2_45_imag;
  wire[46:0] T11207;
  wire[45:0] T11208;
  wire[45:0] T11209;
  wire T11210;
  wire[46:0] T11211;
  wire[46:0] T11212;
  wire T11213;
  wire[46:0] T11214;
  wire[46:0] twiddle4_2_46_imag;
  wire[46:0] T11215;
  wire[45:0] T11216;
  wire[45:0] T11217;
  wire T11218;
  wire[46:0] T11219;
  wire[46:0] T11220;
  wire[46:0] twiddle4_2_47_imag;
  wire[46:0] T11221;
  wire[45:0] T11222;
  wire[45:0] T11223;
  wire T11224;
  wire[46:0] T11225;
  wire[46:0] T11226;
  wire T11227;
  wire T11228;
  wire T11229;
  wire T11230;
  wire[46:0] T11231;
  wire[46:0] T11232;
  wire[46:0] T11233;
  wire[46:0] T11234;
  wire[46:0] twiddle4_2_48_imag;
  wire[46:0] T11235;
  wire[45:0] T11236;
  wire[45:0] T11237;
  wire T11238;
  wire[46:0] T11239;
  wire[46:0] T11240;
  wire[46:0] twiddle4_2_49_imag;
  wire[46:0] T11241;
  wire[45:0] T11242;
  wire[45:0] T11243;
  wire T11244;
  wire[46:0] T11245;
  wire[46:0] T11246;
  wire T11247;
  wire[46:0] T11248;
  wire[46:0] twiddle4_2_50_imag;
  wire[46:0] T11249;
  wire[45:0] T11250;
  wire[45:0] T11251;
  wire T11252;
  wire[46:0] T11253;
  wire[46:0] T11254;
  wire[46:0] twiddle4_2_51_imag;
  wire[46:0] T11255;
  wire[45:0] T11256;
  wire[45:0] T11257;
  wire T11258;
  wire[46:0] T11259;
  wire[46:0] T11260;
  wire T11261;
  wire T11262;
  wire[46:0] T11263;
  wire[46:0] T11264;
  wire[46:0] twiddle4_2_52_imag;
  wire[46:0] T11265;
  wire[45:0] T11266;
  wire[45:0] T11267;
  wire T11268;
  wire[46:0] T11269;
  wire[46:0] T11270;
  wire[46:0] twiddle4_2_53_imag;
  wire[46:0] T11271;
  wire[45:0] T11272;
  wire[45:0] T11273;
  wire T11274;
  wire[46:0] T11275;
  wire[46:0] T11276;
  wire T11277;
  wire[46:0] T11278;
  wire[46:0] twiddle4_2_54_imag;
  wire[46:0] T11279;
  wire[45:0] T11280;
  wire[45:0] T11281;
  wire T11282;
  wire[46:0] T11283;
  wire[46:0] T11284;
  wire[46:0] twiddle4_2_55_imag;
  wire[46:0] T11285;
  wire[45:0] T11286;
  wire[45:0] T11287;
  wire T11288;
  wire[46:0] T11289;
  wire[46:0] T11290;
  wire T11291;
  wire T11292;
  wire T11293;
  wire[46:0] T11294;
  wire[46:0] T11295;
  wire[46:0] T11296;
  wire[46:0] twiddle4_2_56_imag;
  wire[46:0] T11297;
  wire[45:0] T11298;
  wire[45:0] T11299;
  wire T11300;
  wire[46:0] T11301;
  wire[46:0] T11302;
  wire[46:0] twiddle4_2_57_imag;
  wire[46:0] T11303;
  wire[45:0] T11304;
  wire[45:0] T11305;
  wire T11306;
  wire[46:0] T11307;
  wire[46:0] T11308;
  wire T11309;
  wire[46:0] T11310;
  wire[46:0] twiddle4_2_58_imag;
  wire[46:0] T11311;
  wire[45:0] T11312;
  wire[45:0] T11313;
  wire T11314;
  wire[46:0] T11315;
  wire[46:0] T11316;
  wire[46:0] twiddle4_2_59_imag;
  wire[46:0] T11317;
  wire[45:0] T11318;
  wire[45:0] T11319;
  wire T11320;
  wire[46:0] T11321;
  wire[46:0] T11322;
  wire T11323;
  wire T11324;
  wire[46:0] T11325;
  wire[46:0] T11326;
  wire[46:0] twiddle4_2_60_imag;
  wire[46:0] T11327;
  wire[45:0] T11328;
  wire[45:0] T11329;
  wire T11330;
  wire[46:0] T11331;
  wire[46:0] T11332;
  wire[46:0] twiddle4_2_61_imag;
  wire[46:0] T11333;
  wire[45:0] T11334;
  wire[45:0] T11335;
  wire T11336;
  wire[46:0] T11337;
  wire[46:0] T11338;
  wire T11339;
  wire[46:0] T11340;
  wire[46:0] twiddle4_2_62_imag;
  wire[46:0] T11341;
  wire[45:0] T11342;
  wire[45:0] T11343;
  wire T11344;
  wire[46:0] T11345;
  wire[46:0] T11346;
  wire[46:0] twiddle4_2_63_imag;
  wire[46:0] T11347;
  wire[45:0] T11348;
  wire[45:0] T11349;
  wire T11350;
  wire[46:0] T11351;
  wire[46:0] T11352;
  wire T11353;
  wire T11354;
  wire T11355;
  wire T11356;
  wire T11357;
  wire T11358;
  wire T11359;
  wire[47:0] T11360;
  wire[46:0] T11361;
  wire[46:0] T11362;
  wire[46:0] T11363;
  wire[46:0] T11364;
  wire[46:0] T11365;
  wire[46:0] T11366;
  wire[46:0] twiddle4_2_64_imag;
  wire[46:0] T11367;
  wire[45:0] T11368;
  wire[45:0] T11369;
  wire T11370;
  wire[46:0] T11371;
  wire[46:0] T11372;
  wire[46:0] twiddle4_2_65_imag;
  wire[46:0] T11373;
  wire[45:0] T11374;
  wire[45:0] T11375;
  wire T11376;
  wire[46:0] T11377;
  wire[46:0] T11378;
  wire T11379;
  wire[46:0] T11380;
  wire[46:0] twiddle4_2_66_imag;
  wire[46:0] T11381;
  wire[45:0] T11382;
  wire[45:0] T11383;
  wire T11384;
  wire[46:0] T11385;
  wire[46:0] T11386;
  wire[46:0] twiddle4_2_67_imag;
  wire[46:0] T11387;
  wire[45:0] T11388;
  wire[45:0] T11389;
  wire T11390;
  wire[46:0] T11391;
  wire[46:0] T11392;
  wire T11393;
  wire T11394;
  wire[46:0] T11395;
  wire[46:0] T11396;
  wire[46:0] twiddle4_2_68_imag;
  wire[46:0] T11397;
  wire[45:0] T11398;
  wire[45:0] T11399;
  wire T11400;
  wire[46:0] T11401;
  wire[46:0] T11402;
  wire[46:0] twiddle4_2_69_imag;
  wire[46:0] T11403;
  wire[45:0] T11404;
  wire[45:0] T11405;
  wire T11406;
  wire[46:0] T11407;
  wire[46:0] T11408;
  wire T11409;
  wire[46:0] T11410;
  wire[46:0] twiddle4_2_70_imag;
  wire[46:0] T11411;
  wire[45:0] T11412;
  wire[45:0] T11413;
  wire T11414;
  wire[46:0] T11415;
  wire[46:0] T11416;
  wire[46:0] twiddle4_2_71_imag;
  wire[46:0] T11417;
  wire[45:0] T11418;
  wire[45:0] T11419;
  wire T11420;
  wire[46:0] T11421;
  wire[46:0] T11422;
  wire T11423;
  wire T11424;
  wire T11425;
  wire[46:0] T11426;
  wire[46:0] T11427;
  wire[46:0] T11428;
  wire[46:0] twiddle4_2_72_imag;
  wire[46:0] T11429;
  wire[45:0] T11430;
  wire[45:0] T11431;
  wire T11432;
  wire[46:0] T11433;
  wire[46:0] T11434;
  wire[46:0] twiddle4_2_73_imag;
  wire[46:0] T11435;
  wire[45:0] T11436;
  wire[45:0] T11437;
  wire T11438;
  wire[46:0] T11439;
  wire[46:0] T11440;
  wire T11441;
  wire[46:0] T11442;
  wire[46:0] twiddle4_2_74_imag;
  wire[46:0] T11443;
  wire[45:0] T11444;
  wire[45:0] T11445;
  wire T11446;
  wire[46:0] T11447;
  wire[46:0] T11448;
  wire[46:0] twiddle4_2_75_imag;
  wire[46:0] T11449;
  wire[45:0] T11450;
  wire[45:0] T11451;
  wire T11452;
  wire[46:0] T11453;
  wire[46:0] T11454;
  wire T11455;
  wire T11456;
  wire[46:0] T11457;
  wire[46:0] T11458;
  wire[46:0] twiddle4_2_76_imag;
  wire[46:0] T11459;
  wire[45:0] T11460;
  wire[45:0] T11461;
  wire T11462;
  wire[46:0] T11463;
  wire[46:0] T11464;
  wire[46:0] twiddle4_2_77_imag;
  wire[46:0] T11465;
  wire[45:0] T11466;
  wire[45:0] T11467;
  wire T11468;
  wire[46:0] T11469;
  wire[46:0] T11470;
  wire T11471;
  wire[46:0] T11472;
  wire[46:0] twiddle4_2_78_imag;
  wire[46:0] T11473;
  wire[45:0] T11474;
  wire[45:0] T11475;
  wire T11476;
  wire[46:0] T11477;
  wire[46:0] T11478;
  wire[46:0] twiddle4_2_79_imag;
  wire[46:0] T11479;
  wire[45:0] T11480;
  wire[45:0] T11481;
  wire T11482;
  wire[46:0] T11483;
  wire[46:0] T11484;
  wire T11485;
  wire T11486;
  wire T11487;
  wire T11488;
  wire[46:0] T11489;
  wire[46:0] T11490;
  wire[46:0] T11491;
  wire[46:0] T11492;
  wire[46:0] twiddle4_2_80_imag;
  wire[46:0] T11493;
  wire[45:0] T11494;
  wire[45:0] T11495;
  wire T11496;
  wire[46:0] T11497;
  wire[46:0] T11498;
  wire[46:0] twiddle4_2_81_imag;
  wire[46:0] T11499;
  wire[45:0] T11500;
  wire[45:0] T11501;
  wire T11502;
  wire[46:0] T11503;
  wire[46:0] T11504;
  wire T11505;
  wire[46:0] T11506;
  wire[46:0] twiddle4_2_82_imag;
  wire[46:0] T11507;
  wire[45:0] T11508;
  wire[45:0] T11509;
  wire T11510;
  wire[46:0] T11511;
  wire[46:0] T11512;
  wire[46:0] twiddle4_2_83_imag;
  wire[46:0] T11513;
  wire[45:0] T11514;
  wire[45:0] T11515;
  wire T11516;
  wire[46:0] T11517;
  wire[46:0] T11518;
  wire T11519;
  wire T11520;
  wire[46:0] T11521;
  wire[46:0] T11522;
  wire[46:0] twiddle4_2_84_imag;
  wire[46:0] T11523;
  wire[45:0] T11524;
  wire[45:0] T11525;
  wire T11526;
  wire[46:0] T11527;
  wire[46:0] T11528;
  wire[46:0] twiddle4_2_85_imag;
  wire[46:0] T11529;
  wire[45:0] T11530;
  wire[45:0] T11531;
  wire T11532;
  wire[46:0] T11533;
  wire[46:0] T11534;
  wire T11535;
  wire[46:0] T11536;
  wire[46:0] twiddle4_2_86_imag;
  wire[46:0] T11537;
  wire[46:0] T11538;
  wire[46:0] T11539;
  wire[46:0] T11540;
  wire[46:0] twiddle4_2_87_imag;
  wire[46:0] T11541;
  wire[46:0] T11542;
  wire[46:0] T11543;
  wire[46:0] T11544;
  wire T11545;
  wire T11546;
  wire T11547;
  wire[46:0] T11548;
  wire[46:0] T11549;
  wire[46:0] T11550;
  wire[46:0] twiddle4_2_88_imag;
  wire[46:0] T11551;
  wire[46:0] T11552;
  wire[46:0] T11553;
  wire[46:0] T11554;
  wire[46:0] twiddle4_2_89_imag;
  wire[46:0] T11555;
  wire[46:0] T11556;
  wire[46:0] T11557;
  wire[46:0] T11558;
  wire T11559;
  wire[46:0] T11560;
  wire[46:0] twiddle4_2_90_imag;
  wire[46:0] T11561;
  wire[46:0] T11562;
  wire[46:0] T11563;
  wire[46:0] T11564;
  wire[46:0] twiddle4_2_91_imag;
  wire[46:0] T11565;
  wire[46:0] T11566;
  wire[46:0] T11567;
  wire[46:0] T11568;
  wire T11569;
  wire T11570;
  wire[46:0] T11571;
  wire[46:0] T11572;
  wire[46:0] twiddle4_2_92_imag;
  wire[46:0] T11573;
  wire[46:0] T11574;
  wire[46:0] T11575;
  wire[46:0] T11576;
  wire[46:0] twiddle4_2_93_imag;
  wire[46:0] T11577;
  wire[46:0] T11578;
  wire[46:0] T11579;
  wire[46:0] T11580;
  wire T11581;
  wire[46:0] T11582;
  wire[46:0] twiddle4_2_94_imag;
  wire[46:0] T11583;
  wire[46:0] T11584;
  wire[46:0] T11585;
  wire[46:0] T11586;
  wire[46:0] twiddle4_2_95_imag;
  wire[46:0] T11587;
  wire[46:0] T11588;
  wire[46:0] T11589;
  wire[46:0] T11590;
  wire T11591;
  wire T11592;
  wire T11593;
  wire T11594;
  wire T11595;
  wire[46:0] T11596;
  wire[46:0] T11597;
  wire[46:0] T11598;
  wire[46:0] T11599;
  wire[46:0] T11600;
  wire[46:0] twiddle4_2_96_imag;
  wire[46:0] T11601;
  wire[46:0] T11602;
  wire[46:0] T11603;
  wire[46:0] T11604;
  wire[46:0] twiddle4_2_97_imag;
  wire[46:0] T11605;
  wire[46:0] T11606;
  wire[46:0] T11607;
  wire[46:0] T11608;
  wire T11609;
  wire[46:0] T11610;
  wire[46:0] twiddle4_2_98_imag;
  wire[46:0] T11611;
  wire[46:0] T11612;
  wire[46:0] T11613;
  wire[46:0] T11614;
  wire[46:0] twiddle4_2_99_imag;
  wire[46:0] T11615;
  wire[46:0] T11616;
  wire[46:0] T11617;
  wire[46:0] T11618;
  wire T11619;
  wire T11620;
  wire[46:0] T11621;
  wire[46:0] T11622;
  wire[46:0] twiddle4_2_100_imag;
  wire[46:0] T11623;
  wire[46:0] T11624;
  wire[46:0] T11625;
  wire[46:0] T11626;
  wire[46:0] twiddle4_2_101_imag;
  wire[46:0] T11627;
  wire[46:0] T11628;
  wire[46:0] T11629;
  wire[46:0] T11630;
  wire T11631;
  wire[46:0] T11632;
  wire[46:0] twiddle4_2_102_imag;
  wire[46:0] T11633;
  wire[46:0] T11634;
  wire[46:0] T11635;
  wire[46:0] T11636;
  wire[46:0] twiddle4_2_103_imag;
  wire[46:0] T11637;
  wire[46:0] T11638;
  wire[46:0] T11639;
  wire[46:0] T11640;
  wire T11641;
  wire T11642;
  wire T11643;
  wire[46:0] T11644;
  wire[46:0] T11645;
  wire[46:0] T11646;
  wire[46:0] twiddle4_2_104_imag;
  wire[46:0] T11647;
  wire[46:0] T11648;
  wire[46:0] T11649;
  wire[46:0] T11650;
  wire[46:0] twiddle4_2_105_imag;
  wire[46:0] T11651;
  wire[46:0] T11652;
  wire[46:0] T11653;
  wire[46:0] T11654;
  wire T11655;
  wire[46:0] T11656;
  wire[46:0] twiddle4_2_106_imag;
  wire[46:0] T11657;
  wire[46:0] T11658;
  wire[46:0] T11659;
  wire[46:0] T11660;
  wire[46:0] twiddle4_2_107_imag;
  wire[46:0] T11661;
  wire[46:0] T11662;
  wire[46:0] T11663;
  wire[46:0] T11664;
  wire T11665;
  wire T11666;
  wire[46:0] T11667;
  wire[46:0] T11668;
  wire[46:0] twiddle4_2_108_imag;
  wire[46:0] T11669;
  wire[46:0] T11670;
  wire[46:0] T11671;
  wire[46:0] T11672;
  wire[46:0] twiddle4_2_109_imag;
  wire[46:0] T11673;
  wire[46:0] T11674;
  wire[46:0] T11675;
  wire[46:0] T11676;
  wire T11677;
  wire[46:0] T11678;
  wire[46:0] twiddle4_2_110_imag;
  wire[46:0] T11679;
  wire[46:0] T11680;
  wire[46:0] T11681;
  wire[46:0] T11682;
  wire[46:0] twiddle4_2_111_imag;
  wire[46:0] T11683;
  wire[46:0] T11684;
  wire[46:0] T11685;
  wire[46:0] T11686;
  wire T11687;
  wire T11688;
  wire T11689;
  wire T11690;
  wire[46:0] T11691;
  wire[46:0] T11692;
  wire[46:0] T11693;
  wire[46:0] T11694;
  wire[46:0] twiddle4_2_112_imag;
  wire[46:0] T11695;
  wire[46:0] T11696;
  wire[46:0] T11697;
  wire[46:0] T11698;
  wire[46:0] twiddle4_2_113_imag;
  wire[46:0] T11699;
  wire[46:0] T11700;
  wire[46:0] T11701;
  wire[46:0] T11702;
  wire T11703;
  wire[46:0] T11704;
  wire[46:0] twiddle4_2_114_imag;
  wire[46:0] T11705;
  wire[46:0] T11706;
  wire[46:0] T11707;
  wire[46:0] T11708;
  wire[46:0] twiddle4_2_115_imag;
  wire[46:0] T11709;
  wire[46:0] T11710;
  wire[46:0] T11711;
  wire[46:0] T11712;
  wire T11713;
  wire T11714;
  wire[46:0] T11715;
  wire[46:0] T11716;
  wire[46:0] twiddle4_2_116_imag;
  wire[46:0] T11717;
  wire[46:0] T11718;
  wire[46:0] T11719;
  wire[46:0] T11720;
  wire[46:0] twiddle4_2_117_imag;
  wire[46:0] T11721;
  wire[46:0] T11722;
  wire[46:0] T11723;
  wire[46:0] T11724;
  wire T11725;
  wire[46:0] T11726;
  wire[46:0] twiddle4_2_118_imag;
  wire[46:0] T11727;
  wire[46:0] T11728;
  wire[46:0] T11729;
  wire[46:0] T11730;
  wire[46:0] twiddle4_2_119_imag;
  wire[46:0] T11731;
  wire[46:0] T11732;
  wire[46:0] T11733;
  wire[46:0] T11734;
  wire T11735;
  wire T11736;
  wire T11737;
  wire[46:0] T11738;
  wire[46:0] T11739;
  wire[46:0] T11740;
  wire[46:0] twiddle4_2_120_imag;
  wire[46:0] T11741;
  wire[46:0] T11742;
  wire[46:0] T11743;
  wire[46:0] T11744;
  wire[46:0] twiddle4_2_121_imag;
  wire[46:0] T11745;
  wire[46:0] T11746;
  wire[46:0] T11747;
  wire[46:0] T11748;
  wire T11749;
  wire[46:0] T11750;
  wire[46:0] twiddle4_2_122_imag;
  wire[46:0] T11751;
  wire[46:0] T11752;
  wire[46:0] T11753;
  wire[46:0] T11754;
  wire[46:0] twiddle4_2_123_imag;
  wire[46:0] T11755;
  wire[46:0] T11756;
  wire[46:0] T11757;
  wire[46:0] T11758;
  wire T11759;
  wire T11760;
  wire[46:0] T11761;
  wire[46:0] T11762;
  wire[46:0] twiddle4_2_124_imag;
  wire[46:0] T11763;
  wire[46:0] T11764;
  wire[46:0] T11765;
  wire[46:0] T11766;
  wire[46:0] twiddle4_2_125_imag;
  wire[46:0] T11767;
  wire[46:0] T11768;
  wire[46:0] T11769;
  wire[46:0] T11770;
  wire T11771;
  wire[46:0] T11772;
  wire[46:0] twiddle4_2_126_imag;
  wire[46:0] T11773;
  wire[46:0] T11774;
  wire[46:0] T11775;
  wire[46:0] T11776;
  wire[46:0] twiddle4_2_127_imag;
  wire[46:0] T11777;
  wire[46:0] T11778;
  wire[46:0] T11779;
  wire[46:0] T11780;
  wire T11781;
  wire T11782;
  wire T11783;
  wire T11784;
  wire T11785;
  wire T11786;
  wire T11787;
  wire T11788;
  wire[47:0] T11789;
  wire[46:0] T11790;
  wire[46:0] T11791;
  wire[46:0] T11792;
  wire[46:0] T11793;
  wire[46:0] T11794;
  wire[46:0] T11795;
  wire[46:0] T11796;
  wire[46:0] twiddle4_2_128_imag;
  wire[46:0] T11797;
  wire[46:0] T11798;
  wire[46:0] T11799;
  wire[46:0] T11800;
  wire[46:0] twiddle4_2_129_imag;
  wire[46:0] T11801;
  wire[46:0] T11802;
  wire[46:0] T11803;
  wire[46:0] T11804;
  wire T11805;
  wire[46:0] T11806;
  wire[46:0] twiddle4_2_130_imag;
  wire[46:0] T11807;
  wire[46:0] T11808;
  wire[46:0] T11809;
  wire[46:0] T11810;
  wire[46:0] twiddle4_2_131_imag;
  wire[46:0] T11811;
  wire[46:0] T11812;
  wire[46:0] T11813;
  wire[46:0] T11814;
  wire T11815;
  wire T11816;
  wire[46:0] T11817;
  wire[46:0] T11818;
  wire[46:0] twiddle4_2_132_imag;
  wire[46:0] T11819;
  wire[46:0] T11820;
  wire[46:0] T11821;
  wire[46:0] T11822;
  wire[46:0] twiddle4_2_133_imag;
  wire[46:0] T11823;
  wire[46:0] T11824;
  wire[46:0] T11825;
  wire[46:0] T11826;
  wire T11827;
  wire[46:0] T11828;
  wire[46:0] twiddle4_2_134_imag;
  wire[46:0] T11829;
  wire[46:0] T11830;
  wire[46:0] T11831;
  wire[46:0] T11832;
  wire[46:0] twiddle4_2_135_imag;
  wire[46:0] T11833;
  wire[46:0] T11834;
  wire[46:0] T11835;
  wire[46:0] T11836;
  wire T11837;
  wire T11838;
  wire T11839;
  wire[46:0] T11840;
  wire[46:0] T11841;
  wire[46:0] T11842;
  wire[46:0] twiddle4_2_136_imag;
  wire[46:0] T11843;
  wire[46:0] T11844;
  wire[46:0] T11845;
  wire[46:0] T11846;
  wire[46:0] twiddle4_2_137_imag;
  wire[46:0] T11847;
  wire[46:0] T11848;
  wire[46:0] T11849;
  wire[46:0] T11850;
  wire T11851;
  wire[46:0] T11852;
  wire[46:0] twiddle4_2_138_imag;
  wire[46:0] T11853;
  wire[46:0] T11854;
  wire[46:0] T11855;
  wire[46:0] T11856;
  wire[46:0] twiddle4_2_139_imag;
  wire[46:0] T11857;
  wire[46:0] T11858;
  wire[46:0] T11859;
  wire[46:0] T11860;
  wire T11861;
  wire T11862;
  wire[46:0] T11863;
  wire[46:0] T11864;
  wire[46:0] twiddle4_2_140_imag;
  wire[46:0] T11865;
  wire[46:0] T11866;
  wire[46:0] T11867;
  wire[46:0] T11868;
  wire[46:0] twiddle4_2_141_imag;
  wire[46:0] T11869;
  wire[46:0] T11870;
  wire[46:0] T11871;
  wire[46:0] T11872;
  wire T11873;
  wire[46:0] T11874;
  wire[46:0] twiddle4_2_142_imag;
  wire[46:0] T11875;
  wire[46:0] T11876;
  wire[46:0] T11877;
  wire[46:0] T11878;
  wire[46:0] twiddle4_2_143_imag;
  wire[46:0] T11879;
  wire[46:0] T11880;
  wire[46:0] T11881;
  wire[46:0] T11882;
  wire T11883;
  wire T11884;
  wire T11885;
  wire T11886;
  wire[46:0] T11887;
  wire[46:0] T11888;
  wire[46:0] T11889;
  wire[46:0] T11890;
  wire[46:0] twiddle4_2_144_imag;
  wire[46:0] T11891;
  wire[46:0] T11892;
  wire[46:0] T11893;
  wire[46:0] T11894;
  wire[46:0] twiddle4_2_145_imag;
  wire[46:0] T11895;
  wire[46:0] T11896;
  wire[46:0] T11897;
  wire[46:0] T11898;
  wire T11899;
  wire[46:0] T11900;
  wire[46:0] twiddle4_2_146_imag;
  wire[46:0] T11901;
  wire[46:0] T11902;
  wire[46:0] T11903;
  wire[46:0] T11904;
  wire[46:0] twiddle4_2_147_imag;
  wire[46:0] T11905;
  wire[46:0] T11906;
  wire[46:0] T11907;
  wire[46:0] T11908;
  wire T11909;
  wire T11910;
  wire[46:0] T11911;
  wire[46:0] T11912;
  wire[46:0] twiddle4_2_148_imag;
  wire[46:0] T11913;
  wire[46:0] T11914;
  wire[46:0] T11915;
  wire[46:0] T11916;
  wire[46:0] twiddle4_2_149_imag;
  wire[46:0] T11917;
  wire[46:0] T11918;
  wire[46:0] T11919;
  wire[46:0] T11920;
  wire T11921;
  wire[46:0] T11922;
  wire[46:0] twiddle4_2_150_imag;
  wire[46:0] T11923;
  wire[46:0] T11924;
  wire[46:0] T11925;
  wire[46:0] T11926;
  wire[46:0] twiddle4_2_151_imag;
  wire[46:0] T11927;
  wire[46:0] T11928;
  wire[46:0] T11929;
  wire[46:0] T11930;
  wire T11931;
  wire T11932;
  wire T11933;
  wire[46:0] T11934;
  wire[46:0] T11935;
  wire[46:0] T11936;
  wire[46:0] twiddle4_2_152_imag;
  wire[46:0] T11937;
  wire[46:0] T11938;
  wire[46:0] T11939;
  wire[46:0] T11940;
  wire[46:0] twiddle4_2_153_imag;
  wire[46:0] T11941;
  wire[46:0] T11942;
  wire[46:0] T11943;
  wire[46:0] T11944;
  wire T11945;
  wire[46:0] T11946;
  wire[46:0] twiddle4_2_154_imag;
  wire[46:0] T11947;
  wire[46:0] T11948;
  wire[46:0] T11949;
  wire[46:0] T11950;
  wire[46:0] twiddle4_2_155_imag;
  wire[46:0] T11951;
  wire[46:0] T11952;
  wire[46:0] T11953;
  wire[46:0] T11954;
  wire T11955;
  wire T11956;
  wire[46:0] T11957;
  wire[46:0] T11958;
  wire[46:0] twiddle4_2_156_imag;
  wire[46:0] T11959;
  wire[46:0] T11960;
  wire[46:0] T11961;
  wire[46:0] T11962;
  wire[46:0] twiddle4_2_157_imag;
  wire[46:0] T11963;
  wire[46:0] T11964;
  wire[46:0] T11965;
  wire[46:0] T11966;
  wire T11967;
  wire[46:0] T11968;
  wire[46:0] twiddle4_2_158_imag;
  wire[46:0] T11969;
  wire[46:0] T11970;
  wire[46:0] T11971;
  wire[46:0] T11972;
  wire[46:0] twiddle4_2_159_imag;
  wire[46:0] T11973;
  wire[46:0] T11974;
  wire[46:0] T11975;
  wire[46:0] T11976;
  wire T11977;
  wire T11978;
  wire T11979;
  wire T11980;
  wire T11981;
  wire[46:0] T11982;
  wire[46:0] T11983;
  wire[46:0] T11984;
  wire[46:0] T11985;
  wire[46:0] T11986;
  wire[46:0] twiddle4_2_160_imag;
  wire[46:0] T11987;
  wire[46:0] T11988;
  wire[46:0] T11989;
  wire[46:0] T11990;
  wire[46:0] twiddle4_2_161_imag;
  wire[46:0] T11991;
  wire[46:0] T11992;
  wire[46:0] T11993;
  wire[46:0] T11994;
  wire T11995;
  wire[46:0] T11996;
  wire[46:0] twiddle4_2_162_imag;
  wire[46:0] T11997;
  wire[46:0] T11998;
  wire[46:0] T11999;
  wire[46:0] T12000;
  wire[46:0] twiddle4_2_163_imag;
  wire[46:0] T12001;
  wire[46:0] T12002;
  wire[46:0] T12003;
  wire[46:0] T12004;
  wire T12005;
  wire T12006;
  wire[46:0] T12007;
  wire[46:0] T12008;
  wire[46:0] twiddle4_2_164_imag;
  wire[46:0] T12009;
  wire[46:0] T12010;
  wire[46:0] T12011;
  wire[46:0] T12012;
  wire[46:0] twiddle4_2_165_imag;
  wire[46:0] T12013;
  wire[46:0] T12014;
  wire[46:0] T12015;
  wire[46:0] T12016;
  wire T12017;
  wire[46:0] T12018;
  wire[46:0] twiddle4_2_166_imag;
  wire[46:0] T12019;
  wire[46:0] T12020;
  wire[46:0] T12021;
  wire[46:0] T12022;
  wire[46:0] twiddle4_2_167_imag;
  wire[46:0] T12023;
  wire[46:0] T12024;
  wire[46:0] T12025;
  wire[46:0] T12026;
  wire T12027;
  wire T12028;
  wire T12029;
  wire[46:0] T12030;
  wire[46:0] T12031;
  wire[46:0] T12032;
  wire[46:0] twiddle4_2_168_imag;
  wire[46:0] T12033;
  wire[46:0] T12034;
  wire[46:0] T12035;
  wire[46:0] T12036;
  wire[46:0] twiddle4_2_169_imag;
  wire[46:0] T12037;
  wire[46:0] T12038;
  wire[46:0] T12039;
  wire[46:0] T12040;
  wire T12041;
  wire[46:0] T12042;
  wire[46:0] twiddle4_2_170_imag;
  wire[46:0] T12043;
  wire[46:0] T12044;
  wire[46:0] T12045;
  wire[46:0] T12046;
  wire[46:0] twiddle4_2_171_imag;
  wire[46:0] T12047;
  wire[46:0] T12048;
  wire[46:0] T12049;
  wire[45:0] T12050;
  wire[45:0] T12051;
  wire T12052;
  wire T12053;
  wire T12054;
  wire[46:0] T12055;
  wire[46:0] T12056;
  wire[46:0] twiddle4_2_172_imag;
  wire[46:0] T12057;
  wire[46:0] T12058;
  wire[46:0] T12059;
  wire[45:0] T12060;
  wire[45:0] T12061;
  wire T12062;
  wire[46:0] twiddle4_2_173_imag;
  wire[46:0] T12063;
  wire[46:0] T12064;
  wire[46:0] T12065;
  wire[45:0] T12066;
  wire[45:0] T12067;
  wire T12068;
  wire T12069;
  wire[46:0] T12070;
  wire[46:0] twiddle4_2_174_imag;
  wire[46:0] T12071;
  wire[46:0] T12072;
  wire[46:0] T12073;
  wire[45:0] T12074;
  wire[45:0] T12075;
  wire T12076;
  wire[46:0] twiddle4_2_175_imag;
  wire[46:0] T12077;
  wire[46:0] T12078;
  wire[46:0] T12079;
  wire[45:0] T12080;
  wire[45:0] T12081;
  wire T12082;
  wire T12083;
  wire T12084;
  wire T12085;
  wire T12086;
  wire[46:0] T12087;
  wire[46:0] T12088;
  wire[46:0] T12089;
  wire[46:0] T12090;
  wire[46:0] twiddle4_2_176_imag;
  wire[46:0] T12091;
  wire[46:0] T12092;
  wire[46:0] T12093;
  wire[45:0] T12094;
  wire[45:0] T12095;
  wire T12096;
  wire[46:0] twiddle4_2_177_imag;
  wire[46:0] T12097;
  wire[46:0] T12098;
  wire[46:0] T12099;
  wire[45:0] T12100;
  wire[45:0] T12101;
  wire T12102;
  wire T12103;
  wire[46:0] T12104;
  wire[46:0] twiddle4_2_178_imag;
  wire[46:0] T12105;
  wire[46:0] T12106;
  wire[46:0] T12107;
  wire[45:0] T12108;
  wire[45:0] T12109;
  wire T12110;
  wire[46:0] twiddle4_2_179_imag;
  wire[46:0] T12111;
  wire[46:0] T12112;
  wire[46:0] T12113;
  wire[45:0] T12114;
  wire[45:0] T12115;
  wire T12116;
  wire T12117;
  wire T12118;
  wire[46:0] T12119;
  wire[46:0] T12120;
  wire[46:0] twiddle4_2_180_imag;
  wire[46:0] T12121;
  wire[46:0] T12122;
  wire[46:0] T12123;
  wire[45:0] T12124;
  wire[45:0] T12125;
  wire T12126;
  wire[46:0] twiddle4_2_181_imag;
  wire[46:0] T12127;
  wire[46:0] T12128;
  wire[46:0] T12129;
  wire[45:0] T12130;
  wire[45:0] T12131;
  wire T12132;
  wire T12133;
  wire[46:0] T12134;
  wire[46:0] twiddle4_2_182_imag;
  wire[46:0] T12135;
  wire[46:0] T12136;
  wire[46:0] T12137;
  wire[45:0] T12138;
  wire[45:0] T12139;
  wire T12140;
  wire[46:0] twiddle4_2_183_imag;
  wire[46:0] T12141;
  wire[46:0] T12142;
  wire[46:0] T12143;
  wire[45:0] T12144;
  wire[45:0] T12145;
  wire T12146;
  wire T12147;
  wire T12148;
  wire T12149;
  wire[46:0] T12150;
  wire[46:0] T12151;
  wire[46:0] T12152;
  wire[46:0] twiddle4_2_184_imag;
  wire[46:0] T12153;
  wire[46:0] T12154;
  wire[46:0] T12155;
  wire[45:0] T12156;
  wire[45:0] T12157;
  wire T12158;
  wire[46:0] twiddle4_2_185_imag;
  wire[46:0] T12159;
  wire[46:0] T12160;
  wire[46:0] T12161;
  wire[45:0] T12162;
  wire[45:0] T12163;
  wire T12164;
  wire T12165;
  wire[46:0] T12166;
  wire[46:0] twiddle4_2_186_imag;
  wire[46:0] T12167;
  wire[46:0] T12168;
  wire[46:0] T12169;
  wire[45:0] T12170;
  wire[45:0] T12171;
  wire T12172;
  wire[46:0] twiddle4_2_187_imag;
  wire[46:0] T12173;
  wire[46:0] T12174;
  wire[46:0] T12175;
  wire[45:0] T12176;
  wire[45:0] T12177;
  wire T12178;
  wire T12179;
  wire T12180;
  wire[46:0] T12181;
  wire[46:0] T12182;
  wire[46:0] twiddle4_2_188_imag;
  wire[46:0] T12183;
  wire[46:0] T12184;
  wire[46:0] T12185;
  wire[45:0] T12186;
  wire[45:0] T12187;
  wire T12188;
  wire[46:0] twiddle4_2_189_imag;
  wire[46:0] T12189;
  wire[46:0] T12190;
  wire[46:0] T12191;
  wire[45:0] T12192;
  wire[45:0] T12193;
  wire T12194;
  wire T12195;
  wire[46:0] T12196;
  wire[46:0] twiddle4_2_190_imag;
  wire[46:0] T12197;
  wire[46:0] T12198;
  wire[46:0] T12199;
  wire[45:0] T12200;
  wire[45:0] T12201;
  wire T12202;
  wire[46:0] twiddle4_2_191_imag;
  wire[46:0] T12203;
  wire[46:0] T12204;
  wire[46:0] T12205;
  wire[45:0] T12206;
  wire[45:0] T12207;
  wire T12208;
  wire T12209;
  wire T12210;
  wire T12211;
  wire T12212;
  wire T12213;
  wire T12214;
  wire[46:0] T12215;
  wire[46:0] T12216;
  wire[46:0] T12217;
  wire[46:0] T12218;
  wire[46:0] T12219;
  wire[46:0] T12220;
  wire[46:0] twiddle4_2_192_imag;
  wire[46:0] T12221;
  wire[46:0] T12222;
  wire[46:0] T12223;
  wire[45:0] T12224;
  wire[45:0] T12225;
  wire T12226;
  wire[46:0] twiddle4_2_193_imag;
  wire[46:0] T12227;
  wire[46:0] T12228;
  wire[46:0] T12229;
  wire[45:0] T12230;
  wire[45:0] T12231;
  wire T12232;
  wire T12233;
  wire[46:0] T12234;
  wire[46:0] twiddle4_2_194_imag;
  wire[46:0] T12235;
  wire[46:0] T12236;
  wire[46:0] T12237;
  wire[45:0] T12238;
  wire[45:0] T12239;
  wire T12240;
  wire[46:0] twiddle4_2_195_imag;
  wire[46:0] T12241;
  wire[46:0] T12242;
  wire[46:0] T12243;
  wire[45:0] T12244;
  wire[45:0] T12245;
  wire T12246;
  wire T12247;
  wire T12248;
  wire[46:0] T12249;
  wire[46:0] T12250;
  wire[46:0] twiddle4_2_196_imag;
  wire[46:0] T12251;
  wire[46:0] T12252;
  wire[46:0] T12253;
  wire[45:0] T12254;
  wire[45:0] T12255;
  wire T12256;
  wire[46:0] twiddle4_2_197_imag;
  wire[46:0] T12257;
  wire[46:0] T12258;
  wire[46:0] T12259;
  wire[45:0] T12260;
  wire[45:0] T12261;
  wire T12262;
  wire T12263;
  wire[46:0] T12264;
  wire[46:0] twiddle4_2_198_imag;
  wire[46:0] T12265;
  wire[46:0] T12266;
  wire[46:0] T12267;
  wire[45:0] T12268;
  wire[45:0] T12269;
  wire T12270;
  wire[46:0] twiddle4_2_199_imag;
  wire[46:0] T12271;
  wire[46:0] T12272;
  wire[46:0] T12273;
  wire[45:0] T12274;
  wire[45:0] T12275;
  wire T12276;
  wire T12277;
  wire T12278;
  wire T12279;
  wire[46:0] T12280;
  wire[46:0] T12281;
  wire[46:0] T12282;
  wire[46:0] twiddle4_2_200_imag;
  wire[46:0] T12283;
  wire[46:0] T12284;
  wire[46:0] T12285;
  wire[45:0] T12286;
  wire[45:0] T12287;
  wire T12288;
  wire[46:0] twiddle4_2_201_imag;
  wire[46:0] T12289;
  wire[46:0] T12290;
  wire[46:0] T12291;
  wire[45:0] T12292;
  wire[45:0] T12293;
  wire T12294;
  wire T12295;
  wire[46:0] T12296;
  wire[46:0] twiddle4_2_202_imag;
  wire[46:0] T12297;
  wire[46:0] T12298;
  wire[46:0] T12299;
  wire[45:0] T12300;
  wire[45:0] T12301;
  wire T12302;
  wire[46:0] twiddle4_2_203_imag;
  wire[46:0] T12303;
  wire[46:0] T12304;
  wire[46:0] T12305;
  wire[45:0] T12306;
  wire[45:0] T12307;
  wire T12308;
  wire T12309;
  wire T12310;
  wire[46:0] T12311;
  wire[46:0] T12312;
  wire[46:0] twiddle4_2_204_imag;
  wire[46:0] T12313;
  wire[46:0] T12314;
  wire[46:0] T12315;
  wire[45:0] T12316;
  wire[45:0] T12317;
  wire T12318;
  wire[46:0] twiddle4_2_205_imag;
  wire[46:0] T12319;
  wire[46:0] T12320;
  wire[46:0] T12321;
  wire[45:0] T12322;
  wire[45:0] T12323;
  wire T12324;
  wire T12325;
  wire[46:0] T12326;
  wire[46:0] twiddle4_2_206_imag;
  wire[46:0] T12327;
  wire[46:0] T12328;
  wire[46:0] T12329;
  wire[45:0] T12330;
  wire[45:0] T12331;
  wire T12332;
  wire[46:0] twiddle4_2_207_imag;
  wire[46:0] T12333;
  wire[46:0] T12334;
  wire[46:0] T12335;
  wire[45:0] T12336;
  wire[45:0] T12337;
  wire T12338;
  wire T12339;
  wire T12340;
  wire T12341;
  wire T12342;
  wire[46:0] T12343;
  wire[46:0] T12344;
  wire[46:0] T12345;
  wire[46:0] T12346;
  wire[46:0] twiddle4_2_208_imag;
  wire[46:0] T12347;
  wire[46:0] T12348;
  wire[46:0] T12349;
  wire[45:0] T12350;
  wire[45:0] T12351;
  wire T12352;
  wire[46:0] twiddle4_2_209_imag;
  wire[46:0] T12353;
  wire[46:0] T12354;
  wire[46:0] T12355;
  wire[45:0] T12356;
  wire[45:0] T12357;
  wire T12358;
  wire T12359;
  wire[46:0] T12360;
  wire[46:0] twiddle4_2_210_imag;
  wire[46:0] T12361;
  wire[46:0] T12362;
  wire[46:0] T12363;
  wire[45:0] T12364;
  wire[45:0] T12365;
  wire T12366;
  wire[46:0] twiddle4_2_211_imag;
  wire[46:0] T12367;
  wire[46:0] T12368;
  wire[46:0] T12369;
  wire[45:0] T12370;
  wire[45:0] T12371;
  wire T12372;
  wire T12373;
  wire T12374;
  wire[46:0] T12375;
  wire[46:0] T12376;
  wire[46:0] twiddle4_2_212_imag;
  wire[46:0] T12377;
  wire[46:0] T12378;
  wire[46:0] T12379;
  wire[45:0] T12380;
  wire[45:0] T12381;
  wire T12382;
  wire[46:0] twiddle4_2_213_imag;
  wire[46:0] T12383;
  wire[46:0] T12384;
  wire[46:0] T12385;
  wire[45:0] T12386;
  wire[45:0] T12387;
  wire T12388;
  wire T12389;
  wire[46:0] T12390;
  wire[46:0] twiddle4_2_214_imag;
  wire[46:0] T12391;
  wire[46:0] T12392;
  wire[46:0] T12393;
  wire[45:0] T12394;
  wire[45:0] T12395;
  wire T12396;
  wire[46:0] twiddle4_2_215_imag;
  wire[46:0] T12397;
  wire[46:0] T12398;
  wire[46:0] T12399;
  wire[44:0] T12400;
  wire[44:0] T12401;
  wire[1:0] T12402;
  wire T12403;
  wire T12404;
  wire T12405;
  wire T12406;
  wire[46:0] T12407;
  wire[46:0] T12408;
  wire[46:0] T12409;
  wire[46:0] twiddle4_2_216_imag;
  wire[46:0] T12410;
  wire[46:0] T12411;
  wire[46:0] T12412;
  wire[44:0] T12413;
  wire[44:0] T12414;
  wire[1:0] T12415;
  wire T12416;
  wire[46:0] twiddle4_2_217_imag;
  wire[46:0] T12417;
  wire[46:0] T12418;
  wire[46:0] T12419;
  wire[44:0] T12420;
  wire[44:0] T12421;
  wire[1:0] T12422;
  wire T12423;
  wire T12424;
  wire[46:0] T12425;
  wire[46:0] twiddle4_2_218_imag;
  wire[46:0] T12426;
  wire[46:0] T12427;
  wire[46:0] T12428;
  wire[44:0] T12429;
  wire[44:0] T12430;
  wire[1:0] T12431;
  wire T12432;
  wire[46:0] twiddle4_2_219_imag;
  wire[46:0] T12433;
  wire[46:0] T12434;
  wire[46:0] T12435;
  wire[44:0] T12436;
  wire[44:0] T12437;
  wire[1:0] T12438;
  wire T12439;
  wire T12440;
  wire T12441;
  wire[46:0] T12442;
  wire[46:0] T12443;
  wire[46:0] twiddle4_2_220_imag;
  wire[46:0] T12444;
  wire[46:0] T12445;
  wire[46:0] T12446;
  wire[44:0] T12447;
  wire[44:0] T12448;
  wire[1:0] T12449;
  wire T12450;
  wire[46:0] twiddle4_2_221_imag;
  wire[46:0] T12451;
  wire[46:0] T12452;
  wire[46:0] T12453;
  wire[44:0] T12454;
  wire[44:0] T12455;
  wire[1:0] T12456;
  wire T12457;
  wire T12458;
  wire[46:0] T12459;
  wire[46:0] twiddle4_2_222_imag;
  wire[46:0] T12460;
  wire[46:0] T12461;
  wire[46:0] T12462;
  wire[44:0] T12463;
  wire[44:0] T12464;
  wire[1:0] T12465;
  wire T12466;
  wire[46:0] twiddle4_2_223_imag;
  wire[46:0] T12467;
  wire[46:0] T12468;
  wire[46:0] T12469;
  wire[44:0] T12470;
  wire[44:0] T12471;
  wire[1:0] T12472;
  wire T12473;
  wire T12474;
  wire T12475;
  wire T12476;
  wire T12477;
  wire T12478;
  wire[46:0] T12479;
  wire[46:0] T12480;
  wire[46:0] T12481;
  wire[46:0] T12482;
  wire[46:0] T12483;
  wire[46:0] twiddle4_2_224_imag;
  wire[46:0] T12484;
  wire[46:0] T12485;
  wire[46:0] T12486;
  wire[44:0] T12487;
  wire[44:0] T12488;
  wire[1:0] T12489;
  wire T12490;
  wire[46:0] twiddle4_2_225_imag;
  wire[46:0] T12491;
  wire[46:0] T12492;
  wire[46:0] T12493;
  wire[44:0] T12494;
  wire[44:0] T12495;
  wire[1:0] T12496;
  wire T12497;
  wire T12498;
  wire[46:0] T12499;
  wire[46:0] twiddle4_2_226_imag;
  wire[46:0] T12500;
  wire[46:0] T12501;
  wire[46:0] T12502;
  wire[44:0] T12503;
  wire[44:0] T12504;
  wire[1:0] T12505;
  wire T12506;
  wire[46:0] twiddle4_2_227_imag;
  wire[46:0] T12507;
  wire[46:0] T12508;
  wire[46:0] T12509;
  wire[44:0] T12510;
  wire[44:0] T12511;
  wire[1:0] T12512;
  wire T12513;
  wire T12514;
  wire T12515;
  wire[46:0] T12516;
  wire[46:0] T12517;
  wire[46:0] twiddle4_2_228_imag;
  wire[46:0] T12518;
  wire[46:0] T12519;
  wire[46:0] T12520;
  wire[44:0] T12521;
  wire[44:0] T12522;
  wire[1:0] T12523;
  wire T12524;
  wire[46:0] twiddle4_2_229_imag;
  wire[46:0] T12525;
  wire[46:0] T12526;
  wire[46:0] T12527;
  wire[44:0] T12528;
  wire[44:0] T12529;
  wire[1:0] T12530;
  wire T12531;
  wire T12532;
  wire[46:0] T12533;
  wire[46:0] twiddle4_2_230_imag;
  wire[46:0] T12534;
  wire[46:0] T12535;
  wire[46:0] T12536;
  wire[44:0] T12537;
  wire[44:0] T12538;
  wire[1:0] T12539;
  wire T12540;
  wire[46:0] twiddle4_2_231_imag;
  wire[46:0] T12541;
  wire[46:0] T12542;
  wire[46:0] T12543;
  wire[44:0] T12544;
  wire[44:0] T12545;
  wire[1:0] T12546;
  wire T12547;
  wire T12548;
  wire T12549;
  wire T12550;
  wire[46:0] T12551;
  wire[46:0] T12552;
  wire[46:0] T12553;
  wire[46:0] twiddle4_2_232_imag;
  wire[46:0] T12554;
  wire[46:0] T12555;
  wire[46:0] T12556;
  wire[44:0] T12557;
  wire[44:0] T12558;
  wire[1:0] T12559;
  wire T12560;
  wire[46:0] twiddle4_2_233_imag;
  wire[46:0] T12561;
  wire[46:0] T12562;
  wire[46:0] T12563;
  wire[44:0] T12564;
  wire[44:0] T12565;
  wire[1:0] T12566;
  wire T12567;
  wire T12568;
  wire[46:0] T12569;
  wire[46:0] twiddle4_2_234_imag;
  wire[46:0] T12570;
  wire[46:0] T12571;
  wire[46:0] T12572;
  wire[44:0] T12573;
  wire[44:0] T12574;
  wire[1:0] T12575;
  wire T12576;
  wire[46:0] twiddle4_2_235_imag;
  wire[46:0] T12577;
  wire[46:0] T12578;
  wire[46:0] T12579;
  wire[44:0] T12580;
  wire[44:0] T12581;
  wire[1:0] T12582;
  wire T12583;
  wire T12584;
  wire T12585;
  wire[46:0] T12586;
  wire[46:0] T12587;
  wire[46:0] twiddle4_2_236_imag;
  wire[46:0] T12588;
  wire[46:0] T12589;
  wire[46:0] T12590;
  wire[43:0] T12591;
  wire[43:0] T12592;
  wire[2:0] T12593;
  wire T12594;
  wire[46:0] twiddle4_2_237_imag;
  wire[46:0] T12595;
  wire[46:0] T12596;
  wire[46:0] T12597;
  wire[43:0] T12598;
  wire[43:0] T12599;
  wire[2:0] T12600;
  wire T12601;
  wire T12602;
  wire[46:0] T12603;
  wire[46:0] twiddle4_2_238_imag;
  wire[46:0] T12604;
  wire[46:0] T12605;
  wire[46:0] T12606;
  wire[43:0] T12607;
  wire[43:0] T12608;
  wire[2:0] T12609;
  wire T12610;
  wire[46:0] twiddle4_2_239_imag;
  wire[46:0] T12611;
  wire[46:0] T12612;
  wire[46:0] T12613;
  wire[43:0] T12614;
  wire[43:0] T12615;
  wire[2:0] T12616;
  wire T12617;
  wire T12618;
  wire T12619;
  wire T12620;
  wire T12621;
  wire[46:0] T12622;
  wire[46:0] T12623;
  wire[46:0] T12624;
  wire[46:0] T12625;
  wire[46:0] twiddle4_2_240_imag;
  wire[46:0] T12626;
  wire[46:0] T12627;
  wire[46:0] T12628;
  wire[43:0] T12629;
  wire[43:0] T12630;
  wire[2:0] T12631;
  wire T12632;
  wire[46:0] twiddle4_2_241_imag;
  wire[46:0] T12633;
  wire[46:0] T12634;
  wire[46:0] T12635;
  wire[43:0] T12636;
  wire[43:0] T12637;
  wire[2:0] T12638;
  wire T12639;
  wire T12640;
  wire[46:0] T12641;
  wire[46:0] twiddle4_2_242_imag;
  wire[46:0] T12642;
  wire[46:0] T12643;
  wire[46:0] T12644;
  wire[43:0] T12645;
  wire[43:0] T12646;
  wire[2:0] T12647;
  wire T12648;
  wire[46:0] twiddle4_2_243_imag;
  wire[46:0] T12649;
  wire[46:0] T12650;
  wire[46:0] T12651;
  wire[43:0] T12652;
  wire[43:0] T12653;
  wire[2:0] T12654;
  wire T12655;
  wire T12656;
  wire T12657;
  wire[46:0] T12658;
  wire[46:0] T12659;
  wire[46:0] twiddle4_2_244_imag;
  wire[46:0] T12660;
  wire[46:0] T12661;
  wire[46:0] T12662;
  wire[43:0] T12663;
  wire[43:0] T12664;
  wire[2:0] T12665;
  wire T12666;
  wire[46:0] twiddle4_2_245_imag;
  wire[46:0] T12667;
  wire[46:0] T12668;
  wire[46:0] T12669;
  wire[43:0] T12670;
  wire[43:0] T12671;
  wire[2:0] T12672;
  wire T12673;
  wire T12674;
  wire[46:0] T12675;
  wire[46:0] twiddle4_2_246_imag;
  wire[46:0] T12676;
  wire[46:0] T12677;
  wire[46:0] T12678;
  wire[42:0] T12679;
  wire[42:0] T12680;
  wire[3:0] T12681;
  wire T12682;
  wire[46:0] twiddle4_2_247_imag;
  wire[46:0] T12683;
  wire[46:0] T12684;
  wire[46:0] T12685;
  wire[42:0] T12686;
  wire[42:0] T12687;
  wire[3:0] T12688;
  wire T12689;
  wire T12690;
  wire T12691;
  wire T12692;
  wire[46:0] T12693;
  wire[46:0] T12694;
  wire[46:0] T12695;
  wire[46:0] twiddle4_2_248_imag;
  wire[46:0] T12696;
  wire[46:0] T12697;
  wire[46:0] T12698;
  wire[42:0] T12699;
  wire[42:0] T12700;
  wire[3:0] T12701;
  wire T12702;
  wire[46:0] twiddle4_2_249_imag;
  wire[46:0] T12703;
  wire[46:0] T12704;
  wire[46:0] T12705;
  wire[42:0] T12706;
  wire[42:0] T12707;
  wire[3:0] T12708;
  wire T12709;
  wire T12710;
  wire[46:0] T12711;
  wire[46:0] twiddle4_2_250_imag;
  wire[46:0] T12712;
  wire[46:0] T12713;
  wire[46:0] T12714;
  wire[42:0] T12715;
  wire[42:0] T12716;
  wire[3:0] T12717;
  wire T12718;
  wire[46:0] twiddle4_2_251_imag;
  wire[46:0] T12719;
  wire[46:0] T12720;
  wire[46:0] T12721;
  wire[41:0] T12722;
  wire[41:0] T12723;
  wire[4:0] T12724;
  wire T12725;
  wire T12726;
  wire T12727;
  wire[46:0] T12728;
  wire[46:0] T12729;
  wire[46:0] twiddle4_2_252_imag;
  wire[46:0] T12730;
  wire[46:0] T12731;
  wire[46:0] T12732;
  wire[41:0] T12733;
  wire[41:0] T12734;
  wire[4:0] T12735;
  wire T12736;
  wire[46:0] twiddle4_2_253_imag;
  wire[46:0] T12737;
  wire[46:0] T12738;
  wire[46:0] T12739;
  wire[41:0] T12740;
  wire[41:0] T12741;
  wire[4:0] T12742;
  wire T12743;
  wire T12744;
  wire[46:0] T12745;
  wire[46:0] twiddle4_2_254_imag;
  wire[46:0] T12746;
  wire[46:0] T12747;
  wire[46:0] T12748;
  wire[40:0] T12749;
  wire[40:0] T12750;
  wire[5:0] T12751;
  wire T12752;
  wire[46:0] twiddle4_2_255_imag;
  wire[46:0] T12753;
  wire[46:0] T12754;
  wire[46:0] T12755;
  wire[39:0] T12756;
  wire[39:0] T12757;
  wire[6:0] T12758;
  wire T12759;
  wire T12760;
  wire T12761;
  wire T12762;
  wire T12763;
  wire T12764;
  wire T12765;
  wire T12766;
  wire T12767;
  wire T12768;
  wire[47:0] T12769;
  wire[47:0] T12770;
  wire[47:0] T12771;
  wire[47:0] T12772;
  wire[47:0] T12773;
  wire[47:0] T12774;
  wire[47:0] T12775;
  wire[47:0] T12776;
  wire[47:0] twiddle4_2_256_imag;
  wire[47:0] T12777;
  wire[47:0] T12778;
  wire[47:0] T12779;
  wire[16:0] T12780;
  wire[16:0] T12781;
  wire[30:0] T12782;
  wire T12783;
  wire[47:0] T12784;
  wire[46:0] twiddle4_2_257_imag;
  wire[46:0] T12785;
  wire[46:0] T12786;
  wire[46:0] T12787;
  wire[39:0] T12788;
  wire[39:0] T12789;
  wire[6:0] T12790;
  wire T12791;
  wire T12792;
  wire T12793;
  wire[47:0] T12794;
  wire[46:0] T12795;
  wire[46:0] twiddle4_2_258_imag;
  wire[46:0] T12796;
  wire[46:0] T12797;
  wire[46:0] T12798;
  wire[40:0] T12799;
  wire[40:0] T12800;
  wire[5:0] T12801;
  wire T12802;
  wire[46:0] twiddle4_2_259_imag;
  wire[46:0] T12803;
  wire[46:0] T12804;
  wire[46:0] T12805;
  wire[41:0] T12806;
  wire[41:0] T12807;
  wire[4:0] T12808;
  wire T12809;
  wire T12810;
  wire T12811;
  wire T12812;
  wire[47:0] T12813;
  wire[46:0] T12814;
  wire[46:0] T12815;
  wire[46:0] twiddle4_2_260_imag;
  wire[46:0] T12816;
  wire[46:0] T12817;
  wire[46:0] T12818;
  wire[41:0] T12819;
  wire[41:0] T12820;
  wire[4:0] T12821;
  wire T12822;
  wire[46:0] twiddle4_2_261_imag;
  wire[46:0] T12823;
  wire[46:0] T12824;
  wire[46:0] T12825;
  wire[41:0] T12826;
  wire[41:0] T12827;
  wire[4:0] T12828;
  wire T12829;
  wire T12830;
  wire[46:0] T12831;
  wire[46:0] twiddle4_2_262_imag;
  wire[46:0] T12832;
  wire[46:0] T12833;
  wire[46:0] T12834;
  wire[42:0] T12835;
  wire[42:0] T12836;
  wire[3:0] T12837;
  wire T12838;
  wire[46:0] twiddle4_2_263_imag;
  wire[46:0] T12839;
  wire[46:0] T12840;
  wire[46:0] T12841;
  wire[42:0] T12842;
  wire[42:0] T12843;
  wire[3:0] T12844;
  wire T12845;
  wire T12846;
  wire T12847;
  wire T12848;
  wire T12849;
  wire[47:0] T12850;
  wire[46:0] T12851;
  wire[46:0] T12852;
  wire[46:0] T12853;
  wire[46:0] twiddle4_2_264_imag;
  wire[46:0] T12854;
  wire[46:0] T12855;
  wire[46:0] T12856;
  wire[42:0] T12857;
  wire[42:0] T12858;
  wire[3:0] T12859;
  wire T12860;
  wire[46:0] twiddle4_2_265_imag;
  wire[46:0] T12861;
  wire[46:0] T12862;
  wire[46:0] T12863;
  wire[42:0] T12864;
  wire[42:0] T12865;
  wire[3:0] T12866;
  wire T12867;
  wire T12868;
  wire[46:0] T12869;
  wire[46:0] twiddle4_2_266_imag;
  wire[46:0] T12870;
  wire[46:0] T12871;
  wire[46:0] T12872;
  wire[42:0] T12873;
  wire[42:0] T12874;
  wire[3:0] T12875;
  wire T12876;
  wire[46:0] twiddle4_2_267_imag;
  wire[46:0] T12877;
  wire[46:0] T12878;
  wire[46:0] T12879;
  wire[43:0] T12880;
  wire[43:0] T12881;
  wire[2:0] T12882;
  wire T12883;
  wire T12884;
  wire T12885;
  wire[46:0] T12886;
  wire[46:0] T12887;
  wire[46:0] twiddle4_2_268_imag;
  wire[46:0] T12888;
  wire[46:0] T12889;
  wire[46:0] T12890;
  wire[43:0] T12891;
  wire[43:0] T12892;
  wire[2:0] T12893;
  wire T12894;
  wire[46:0] twiddle4_2_269_imag;
  wire[46:0] T12895;
  wire[46:0] T12896;
  wire[46:0] T12897;
  wire[43:0] T12898;
  wire[43:0] T12899;
  wire[2:0] T12900;
  wire T12901;
  wire T12902;
  wire[46:0] T12903;
  wire[46:0] twiddle4_2_270_imag;
  wire[46:0] T12904;
  wire[46:0] T12905;
  wire[46:0] T12906;
  wire[43:0] T12907;
  wire[43:0] T12908;
  wire[2:0] T12909;
  wire T12910;
  wire[46:0] twiddle4_2_271_imag;
  wire[46:0] T12911;
  wire[46:0] T12912;
  wire[46:0] T12913;
  wire[43:0] T12914;
  wire[43:0] T12915;
  wire[2:0] T12916;
  wire T12917;
  wire T12918;
  wire T12919;
  wire T12920;
  wire T12921;
  wire T12922;
  wire[47:0] T12923;
  wire[46:0] T12924;
  wire[46:0] T12925;
  wire[46:0] T12926;
  wire[46:0] T12927;
  wire[46:0] twiddle4_2_272_imag;
  wire[46:0] T12928;
  wire[46:0] T12929;
  wire[46:0] T12930;
  wire[43:0] T12931;
  wire[43:0] T12932;
  wire[2:0] T12933;
  wire T12934;
  wire[46:0] twiddle4_2_273_imag;
  wire[46:0] T12935;
  wire[46:0] T12936;
  wire[46:0] T12937;
  wire[43:0] T12938;
  wire[43:0] T12939;
  wire[2:0] T12940;
  wire T12941;
  wire T12942;
  wire[46:0] T12943;
  wire[46:0] twiddle4_2_274_imag;
  wire[46:0] T12944;
  wire[46:0] T12945;
  wire[46:0] T12946;
  wire[43:0] T12947;
  wire[43:0] T12948;
  wire[2:0] T12949;
  wire T12950;
  wire[46:0] twiddle4_2_275_imag;
  wire[46:0] T12951;
  wire[46:0] T12952;
  wire[46:0] T12953;
  wire[43:0] T12954;
  wire[43:0] T12955;
  wire[2:0] T12956;
  wire T12957;
  wire T12958;
  wire T12959;
  wire[46:0] T12960;
  wire[46:0] T12961;
  wire[46:0] twiddle4_2_276_imag;
  wire[46:0] T12962;
  wire[46:0] T12963;
  wire[46:0] T12964;
  wire[43:0] T12965;
  wire[43:0] T12966;
  wire[2:0] T12967;
  wire T12968;
  wire[46:0] twiddle4_2_277_imag;
  wire[46:0] T12969;
  wire[46:0] T12970;
  wire[46:0] T12971;
  wire[44:0] T12972;
  wire[44:0] T12973;
  wire[1:0] T12974;
  wire T12975;
  wire T12976;
  wire[46:0] T12977;
  wire[46:0] twiddle4_2_278_imag;
  wire[46:0] T12978;
  wire[46:0] T12979;
  wire[46:0] T12980;
  wire[44:0] T12981;
  wire[44:0] T12982;
  wire[1:0] T12983;
  wire T12984;
  wire[46:0] twiddle4_2_279_imag;
  wire[46:0] T12985;
  wire[46:0] T12986;
  wire[46:0] T12987;
  wire[44:0] T12988;
  wire[44:0] T12989;
  wire[1:0] T12990;
  wire T12991;
  wire T12992;
  wire T12993;
  wire T12994;
  wire[46:0] T12995;
  wire[46:0] T12996;
  wire[46:0] T12997;
  wire[46:0] twiddle4_2_280_imag;
  wire[46:0] T12998;
  wire[46:0] T12999;
  wire[46:0] T13000;
  wire[44:0] T13001;
  wire[44:0] T13002;
  wire[1:0] T13003;
  wire T13004;
  wire[46:0] twiddle4_2_281_imag;
  wire[46:0] T13005;
  wire[46:0] T13006;
  wire[46:0] T13007;
  wire[44:0] T13008;
  wire[44:0] T13009;
  wire[1:0] T13010;
  wire T13011;
  wire T13012;
  wire[46:0] T13013;
  wire[46:0] twiddle4_2_282_imag;
  wire[46:0] T13014;
  wire[46:0] T13015;
  wire[46:0] T13016;
  wire[44:0] T13017;
  wire[44:0] T13018;
  wire[1:0] T13019;
  wire T13020;
  wire[46:0] twiddle4_2_283_imag;
  wire[46:0] T13021;
  wire[46:0] T13022;
  wire[46:0] T13023;
  wire[44:0] T13024;
  wire[44:0] T13025;
  wire[1:0] T13026;
  wire T13027;
  wire T13028;
  wire T13029;
  wire[46:0] T13030;
  wire[46:0] T13031;
  wire[46:0] twiddle4_2_284_imag;
  wire[46:0] T13032;
  wire[46:0] T13033;
  wire[46:0] T13034;
  wire[44:0] T13035;
  wire[44:0] T13036;
  wire[1:0] T13037;
  wire T13038;
  wire[46:0] twiddle4_2_285_imag;
  wire[46:0] T13039;
  wire[46:0] T13040;
  wire[46:0] T13041;
  wire[44:0] T13042;
  wire[44:0] T13043;
  wire[1:0] T13044;
  wire T13045;
  wire T13046;
  wire[46:0] T13047;
  wire[46:0] twiddle4_2_286_imag;
  wire[46:0] T13048;
  wire[46:0] T13049;
  wire[46:0] T13050;
  wire[44:0] T13051;
  wire[44:0] T13052;
  wire[1:0] T13053;
  wire T13054;
  wire[46:0] twiddle4_2_287_imag;
  wire[46:0] T13055;
  wire[46:0] T13056;
  wire[46:0] T13057;
  wire[44:0] T13058;
  wire[44:0] T13059;
  wire[1:0] T13060;
  wire T13061;
  wire T13062;
  wire T13063;
  wire T13064;
  wire T13065;
  wire T13066;
  wire T13067;
  wire[47:0] T13068;
  wire[46:0] T13069;
  wire[46:0] T13070;
  wire[46:0] T13071;
  wire[46:0] T13072;
  wire[46:0] T13073;
  wire[46:0] twiddle4_2_288_imag;
  wire[46:0] T13074;
  wire[46:0] T13075;
  wire[46:0] T13076;
  wire[44:0] T13077;
  wire[44:0] T13078;
  wire[1:0] T13079;
  wire T13080;
  wire[46:0] twiddle4_2_289_imag;
  wire[46:0] T13081;
  wire[46:0] T13082;
  wire[46:0] T13083;
  wire[44:0] T13084;
  wire[44:0] T13085;
  wire[1:0] T13086;
  wire T13087;
  wire T13088;
  wire[46:0] T13089;
  wire[46:0] twiddle4_2_290_imag;
  wire[46:0] T13090;
  wire[46:0] T13091;
  wire[46:0] T13092;
  wire[44:0] T13093;
  wire[44:0] T13094;
  wire[1:0] T13095;
  wire T13096;
  wire[46:0] twiddle4_2_291_imag;
  wire[46:0] T13097;
  wire[46:0] T13098;
  wire[46:0] T13099;
  wire[44:0] T13100;
  wire[44:0] T13101;
  wire[1:0] T13102;
  wire T13103;
  wire T13104;
  wire T13105;
  wire[46:0] T13106;
  wire[46:0] T13107;
  wire[46:0] twiddle4_2_292_imag;
  wire[46:0] T13108;
  wire[46:0] T13109;
  wire[46:0] T13110;
  wire[44:0] T13111;
  wire[44:0] T13112;
  wire[1:0] T13113;
  wire T13114;
  wire[46:0] twiddle4_2_293_imag;
  wire[46:0] T13115;
  wire[46:0] T13116;
  wire[46:0] T13117;
  wire[44:0] T13118;
  wire[44:0] T13119;
  wire[1:0] T13120;
  wire T13121;
  wire T13122;
  wire[46:0] T13123;
  wire[46:0] twiddle4_2_294_imag;
  wire[46:0] T13124;
  wire[46:0] T13125;
  wire[46:0] T13126;
  wire[44:0] T13127;
  wire[44:0] T13128;
  wire[1:0] T13129;
  wire T13130;
  wire[46:0] twiddle4_2_295_imag;
  wire[46:0] T13131;
  wire[46:0] T13132;
  wire[46:0] T13133;
  wire[44:0] T13134;
  wire[44:0] T13135;
  wire[1:0] T13136;
  wire T13137;
  wire T13138;
  wire T13139;
  wire T13140;
  wire[46:0] T13141;
  wire[46:0] T13142;
  wire[46:0] T13143;
  wire[46:0] twiddle4_2_296_imag;
  wire[46:0] T13144;
  wire[46:0] T13145;
  wire[46:0] T13146;
  wire[44:0] T13147;
  wire[44:0] T13148;
  wire[1:0] T13149;
  wire T13150;
  wire[46:0] twiddle4_2_297_imag;
  wire[46:0] T13151;
  wire[46:0] T13152;
  wire[46:0] T13153;
  wire[44:0] T13154;
  wire[44:0] T13155;
  wire[1:0] T13156;
  wire T13157;
  wire T13158;
  wire[46:0] T13159;
  wire[46:0] twiddle4_2_298_imag;
  wire[46:0] T13160;
  wire[46:0] T13161;
  wire[46:0] T13162;
  wire[45:0] T13163;
  wire[45:0] T13164;
  wire T13165;
  wire[46:0] twiddle4_2_299_imag;
  wire[46:0] T13166;
  wire[46:0] T13167;
  wire[46:0] T13168;
  wire[45:0] T13169;
  wire[45:0] T13170;
  wire T13171;
  wire T13172;
  wire T13173;
  wire[46:0] T13174;
  wire[46:0] T13175;
  wire[46:0] twiddle4_2_300_imag;
  wire[46:0] T13176;
  wire[46:0] T13177;
  wire[46:0] T13178;
  wire[45:0] T13179;
  wire[45:0] T13180;
  wire T13181;
  wire[46:0] twiddle4_2_301_imag;
  wire[46:0] T13182;
  wire[46:0] T13183;
  wire[46:0] T13184;
  wire[45:0] T13185;
  wire[45:0] T13186;
  wire T13187;
  wire T13188;
  wire[46:0] T13189;
  wire[46:0] twiddle4_2_302_imag;
  wire[46:0] T13190;
  wire[46:0] T13191;
  wire[46:0] T13192;
  wire[45:0] T13193;
  wire[45:0] T13194;
  wire T13195;
  wire[46:0] twiddle4_2_303_imag;
  wire[46:0] T13196;
  wire[46:0] T13197;
  wire[46:0] T13198;
  wire[45:0] T13199;
  wire[45:0] T13200;
  wire T13201;
  wire T13202;
  wire T13203;
  wire T13204;
  wire T13205;
  wire[46:0] T13206;
  wire[46:0] T13207;
  wire[46:0] T13208;
  wire[46:0] T13209;
  wire[46:0] twiddle4_2_304_imag;
  wire[46:0] T13210;
  wire[46:0] T13211;
  wire[46:0] T13212;
  wire[45:0] T13213;
  wire[45:0] T13214;
  wire T13215;
  wire[46:0] twiddle4_2_305_imag;
  wire[46:0] T13216;
  wire[46:0] T13217;
  wire[46:0] T13218;
  wire[45:0] T13219;
  wire[45:0] T13220;
  wire T13221;
  wire T13222;
  wire[46:0] T13223;
  wire[46:0] twiddle4_2_306_imag;
  wire[46:0] T13224;
  wire[46:0] T13225;
  wire[46:0] T13226;
  wire[45:0] T13227;
  wire[45:0] T13228;
  wire T13229;
  wire[46:0] twiddle4_2_307_imag;
  wire[46:0] T13230;
  wire[46:0] T13231;
  wire[46:0] T13232;
  wire[45:0] T13233;
  wire[45:0] T13234;
  wire T13235;
  wire T13236;
  wire T13237;
  wire[46:0] T13238;
  wire[46:0] T13239;
  wire[46:0] twiddle4_2_308_imag;
  wire[46:0] T13240;
  wire[46:0] T13241;
  wire[46:0] T13242;
  wire[45:0] T13243;
  wire[45:0] T13244;
  wire T13245;
  wire[46:0] twiddle4_2_309_imag;
  wire[46:0] T13246;
  wire[46:0] T13247;
  wire[46:0] T13248;
  wire[45:0] T13249;
  wire[45:0] T13250;
  wire T13251;
  wire T13252;
  wire[46:0] T13253;
  wire[46:0] twiddle4_2_310_imag;
  wire[46:0] T13254;
  wire[46:0] T13255;
  wire[46:0] T13256;
  wire[45:0] T13257;
  wire[45:0] T13258;
  wire T13259;
  wire[46:0] twiddle4_2_311_imag;
  wire[46:0] T13260;
  wire[46:0] T13261;
  wire[46:0] T13262;
  wire[45:0] T13263;
  wire[45:0] T13264;
  wire T13265;
  wire T13266;
  wire T13267;
  wire T13268;
  wire[46:0] T13269;
  wire[46:0] T13270;
  wire[46:0] T13271;
  wire[46:0] twiddle4_2_312_imag;
  wire[46:0] T13272;
  wire[46:0] T13273;
  wire[46:0] T13274;
  wire[45:0] T13275;
  wire[45:0] T13276;
  wire T13277;
  wire[46:0] twiddle4_2_313_imag;
  wire[46:0] T13278;
  wire[46:0] T13279;
  wire[46:0] T13280;
  wire[45:0] T13281;
  wire[45:0] T13282;
  wire T13283;
  wire T13284;
  wire[46:0] T13285;
  wire[46:0] twiddle4_2_314_imag;
  wire[46:0] T13286;
  wire[46:0] T13287;
  wire[46:0] T13288;
  wire[45:0] T13289;
  wire[45:0] T13290;
  wire T13291;
  wire[46:0] twiddle4_2_315_imag;
  wire[46:0] T13292;
  wire[46:0] T13293;
  wire[46:0] T13294;
  wire[45:0] T13295;
  wire[45:0] T13296;
  wire T13297;
  wire T13298;
  wire T13299;
  wire[46:0] T13300;
  wire[46:0] T13301;
  wire[46:0] twiddle4_2_316_imag;
  wire[46:0] T13302;
  wire[46:0] T13303;
  wire[46:0] T13304;
  wire[45:0] T13305;
  wire[45:0] T13306;
  wire T13307;
  wire[46:0] twiddle4_2_317_imag;
  wire[46:0] T13308;
  wire[46:0] T13309;
  wire[46:0] T13310;
  wire[45:0] T13311;
  wire[45:0] T13312;
  wire T13313;
  wire T13314;
  wire[46:0] T13315;
  wire[46:0] twiddle4_2_318_imag;
  wire[46:0] T13316;
  wire[46:0] T13317;
  wire[46:0] T13318;
  wire[45:0] T13319;
  wire[45:0] T13320;
  wire T13321;
  wire[46:0] twiddle4_2_319_imag;
  wire[46:0] T13322;
  wire[46:0] T13323;
  wire[46:0] T13324;
  wire[45:0] T13325;
  wire[45:0] T13326;
  wire T13327;
  wire T13328;
  wire T13329;
  wire T13330;
  wire T13331;
  wire T13332;
  wire T13333;
  wire T13334;
  wire[47:0] T13335;
  wire[46:0] T13336;
  wire[46:0] T13337;
  wire[46:0] T13338;
  wire[46:0] T13339;
  wire[46:0] T13340;
  wire[46:0] T13341;
  wire[46:0] twiddle4_2_320_imag;
  wire[46:0] T13342;
  wire[46:0] T13343;
  wire[46:0] T13344;
  wire[45:0] T13345;
  wire[45:0] T13346;
  wire T13347;
  wire[46:0] twiddle4_2_321_imag;
  wire[46:0] T13348;
  wire[46:0] T13349;
  wire[46:0] T13350;
  wire[45:0] T13351;
  wire[45:0] T13352;
  wire T13353;
  wire T13354;
  wire[46:0] T13355;
  wire[46:0] twiddle4_2_322_imag;
  wire[46:0] T13356;
  wire[46:0] T13357;
  wire[46:0] T13358;
  wire[45:0] T13359;
  wire[45:0] T13360;
  wire T13361;
  wire[46:0] twiddle4_2_323_imag;
  wire[46:0] T13362;
  wire[46:0] T13363;
  wire[46:0] T13364;
  wire[45:0] T13365;
  wire[45:0] T13366;
  wire T13367;
  wire T13368;
  wire T13369;
  wire[46:0] T13370;
  wire[46:0] T13371;
  wire[46:0] twiddle4_2_324_imag;
  wire[46:0] T13372;
  wire[46:0] T13373;
  wire[46:0] T13374;
  wire[45:0] T13375;
  wire[45:0] T13376;
  wire T13377;
  wire[46:0] twiddle4_2_325_imag;
  wire[46:0] T13378;
  wire[46:0] T13379;
  wire[46:0] T13380;
  wire[45:0] T13381;
  wire[45:0] T13382;
  wire T13383;
  wire T13384;
  wire[46:0] T13385;
  wire[46:0] twiddle4_2_326_imag;
  wire[46:0] T13386;
  wire[46:0] T13387;
  wire[46:0] T13388;
  wire[45:0] T13389;
  wire[45:0] T13390;
  wire T13391;
  wire[46:0] twiddle4_2_327_imag;
  wire[46:0] T13392;
  wire[46:0] T13393;
  wire[46:0] T13394;
  wire[45:0] T13395;
  wire[45:0] T13396;
  wire T13397;
  wire T13398;
  wire T13399;
  wire T13400;
  wire[46:0] T13401;
  wire[46:0] T13402;
  wire[46:0] T13403;
  wire[46:0] twiddle4_2_328_imag;
  wire[46:0] T13404;
  wire[46:0] T13405;
  wire[46:0] T13406;
  wire[45:0] T13407;
  wire[45:0] T13408;
  wire T13409;
  wire[46:0] twiddle4_2_329_imag;
  wire[46:0] T13410;
  wire[46:0] T13411;
  wire[46:0] T13412;
  wire[45:0] T13413;
  wire[45:0] T13414;
  wire T13415;
  wire T13416;
  wire[46:0] T13417;
  wire[46:0] twiddle4_2_330_imag;
  wire[46:0] T13418;
  wire[46:0] T13419;
  wire[46:0] T13420;
  wire[45:0] T13421;
  wire[45:0] T13422;
  wire T13423;
  wire[46:0] twiddle4_2_331_imag;
  wire[46:0] T13424;
  wire[46:0] T13425;
  wire[46:0] T13426;
  wire[45:0] T13427;
  wire[45:0] T13428;
  wire T13429;
  wire T13430;
  wire T13431;
  wire[46:0] T13432;
  wire[46:0] T13433;
  wire[46:0] twiddle4_2_332_imag;
  wire[46:0] T13434;
  wire[46:0] T13435;
  wire[46:0] T13436;
  wire[45:0] T13437;
  wire[45:0] T13438;
  wire T13439;
  wire[46:0] twiddle4_2_333_imag;
  wire[46:0] T13440;
  wire[46:0] T13441;
  wire[46:0] T13442;
  wire[45:0] T13443;
  wire[45:0] T13444;
  wire T13445;
  wire T13446;
  wire[46:0] T13447;
  wire[46:0] twiddle4_2_334_imag;
  wire[46:0] T13448;
  wire[46:0] T13449;
  wire[46:0] T13450;
  wire[45:0] T13451;
  wire[45:0] T13452;
  wire T13453;
  wire[46:0] twiddle4_2_335_imag;
  wire[46:0] T13454;
  wire[46:0] T13455;
  wire[46:0] T13456;
  wire[45:0] T13457;
  wire[45:0] T13458;
  wire T13459;
  wire T13460;
  wire T13461;
  wire T13462;
  wire T13463;
  wire[46:0] T13464;
  wire[46:0] T13465;
  wire[46:0] T13466;
  wire[46:0] T13467;
  wire[46:0] twiddle4_2_336_imag;
  wire[46:0] T13468;
  wire[46:0] T13469;
  wire[46:0] T13470;
  wire[45:0] T13471;
  wire[45:0] T13472;
  wire T13473;
  wire[46:0] twiddle4_2_337_imag;
  wire[46:0] T13474;
  wire[46:0] T13475;
  wire[46:0] T13476;
  wire[45:0] T13477;
  wire[45:0] T13478;
  wire T13479;
  wire T13480;
  wire[46:0] T13481;
  wire[46:0] twiddle4_2_338_imag;
  wire[46:0] T13482;
  wire[46:0] T13483;
  wire[46:0] T13484;
  wire[45:0] T13485;
  wire[45:0] T13486;
  wire T13487;
  wire[46:0] twiddle4_2_339_imag;
  wire[46:0] T13488;
  wire[46:0] T13489;
  wire[46:0] T13490;
  wire[45:0] T13491;
  wire[45:0] T13492;
  wire T13493;
  wire T13494;
  wire T13495;
  wire[46:0] T13496;
  wire[46:0] T13497;
  wire[46:0] twiddle4_2_340_imag;
  wire[46:0] T13498;
  wire[46:0] T13499;
  wire[46:0] T13500;
  wire[45:0] T13501;
  wire[45:0] T13502;
  wire T13503;
  wire[46:0] twiddle4_2_341_imag;
  wire[46:0] T13504;
  wire[46:0] T13505;
  wire[46:0] T13506;
  wire[45:0] T13507;
  wire[45:0] T13508;
  wire T13509;
  wire T13510;
  wire[46:0] T13511;
  wire[46:0] twiddle4_2_342_imag;
  wire[46:0] T13512;
  wire[46:0] T13513;
  wire[46:0] T13514;
  wire[46:0] T13515;
  wire[46:0] twiddle4_2_343_imag;
  wire[46:0] T13516;
  wire[46:0] T13517;
  wire[46:0] T13518;
  wire[46:0] T13519;
  wire T13520;
  wire T13521;
  wire T13522;
  wire[46:0] T13523;
  wire[46:0] T13524;
  wire[46:0] T13525;
  wire[46:0] twiddle4_2_344_imag;
  wire[46:0] T13526;
  wire[46:0] T13527;
  wire[46:0] T13528;
  wire[46:0] T13529;
  wire[46:0] twiddle4_2_345_imag;
  wire[46:0] T13530;
  wire[46:0] T13531;
  wire[46:0] T13532;
  wire[46:0] T13533;
  wire T13534;
  wire[46:0] T13535;
  wire[46:0] twiddle4_2_346_imag;
  wire[46:0] T13536;
  wire[46:0] T13537;
  wire[46:0] T13538;
  wire[46:0] T13539;
  wire[46:0] twiddle4_2_347_imag;
  wire[46:0] T13540;
  wire[46:0] T13541;
  wire[46:0] T13542;
  wire[46:0] T13543;
  wire T13544;
  wire T13545;
  wire[46:0] T13546;
  wire[46:0] T13547;
  wire[46:0] twiddle4_2_348_imag;
  wire[46:0] T13548;
  wire[46:0] T13549;
  wire[46:0] T13550;
  wire[46:0] T13551;
  wire[46:0] twiddle4_2_349_imag;
  wire[46:0] T13552;
  wire[46:0] T13553;
  wire[46:0] T13554;
  wire[46:0] T13555;
  wire T13556;
  wire[46:0] T13557;
  wire[46:0] twiddle4_2_350_imag;
  wire[46:0] T13558;
  wire[46:0] T13559;
  wire[46:0] T13560;
  wire[46:0] T13561;
  wire[46:0] twiddle4_2_351_imag;
  wire[46:0] T13562;
  wire[46:0] T13563;
  wire[46:0] T13564;
  wire[46:0] T13565;
  wire T13566;
  wire T13567;
  wire T13568;
  wire T13569;
  wire T13570;
  wire[46:0] T13571;
  wire[46:0] T13572;
  wire[46:0] T13573;
  wire[46:0] T13574;
  wire[46:0] T13575;
  wire[46:0] twiddle4_2_352_imag;
  wire[46:0] T13576;
  wire[46:0] T13577;
  wire[46:0] T13578;
  wire[46:0] T13579;
  wire[46:0] twiddle4_2_353_imag;
  wire[46:0] T13580;
  wire[46:0] T13581;
  wire[46:0] T13582;
  wire[46:0] T13583;
  wire T13584;
  wire[46:0] T13585;
  wire[46:0] twiddle4_2_354_imag;
  wire[46:0] T13586;
  wire[46:0] T13587;
  wire[46:0] T13588;
  wire[46:0] T13589;
  wire[46:0] twiddle4_2_355_imag;
  wire[46:0] T13590;
  wire[46:0] T13591;
  wire[46:0] T13592;
  wire[46:0] T13593;
  wire T13594;
  wire T13595;
  wire[46:0] T13596;
  wire[46:0] T13597;
  wire[46:0] twiddle4_2_356_imag;
  wire[46:0] T13598;
  wire[46:0] T13599;
  wire[46:0] T13600;
  wire[46:0] T13601;
  wire[46:0] twiddle4_2_357_imag;
  wire[46:0] T13602;
  wire[46:0] T13603;
  wire[46:0] T13604;
  wire[46:0] T13605;
  wire T13606;
  wire[46:0] T13607;
  wire[46:0] twiddle4_2_358_imag;
  wire[46:0] T13608;
  wire[46:0] T13609;
  wire[46:0] T13610;
  wire[46:0] T13611;
  wire[46:0] twiddle4_2_359_imag;
  wire[46:0] T13612;
  wire[46:0] T13613;
  wire[46:0] T13614;
  wire[46:0] T13615;
  wire T13616;
  wire T13617;
  wire T13618;
  wire[46:0] T13619;
  wire[46:0] T13620;
  wire[46:0] T13621;
  wire[46:0] twiddle4_2_360_imag;
  wire[46:0] T13622;
  wire[46:0] T13623;
  wire[46:0] T13624;
  wire[46:0] T13625;
  wire[46:0] twiddle4_2_361_imag;
  wire[46:0] T13626;
  wire[46:0] T13627;
  wire[46:0] T13628;
  wire[46:0] T13629;
  wire T13630;
  wire[46:0] T13631;
  wire[46:0] twiddle4_2_362_imag;
  wire[46:0] T13632;
  wire[46:0] T13633;
  wire[46:0] T13634;
  wire[46:0] T13635;
  wire[46:0] twiddle4_2_363_imag;
  wire[46:0] T13636;
  wire[46:0] T13637;
  wire[46:0] T13638;
  wire[46:0] T13639;
  wire T13640;
  wire T13641;
  wire[46:0] T13642;
  wire[46:0] T13643;
  wire[46:0] twiddle4_2_364_imag;
  wire[46:0] T13644;
  wire[46:0] T13645;
  wire[46:0] T13646;
  wire[46:0] T13647;
  wire[46:0] twiddle4_2_365_imag;
  wire[46:0] T13648;
  wire[46:0] T13649;
  wire[46:0] T13650;
  wire[46:0] T13651;
  wire T13652;
  wire[46:0] T13653;
  wire[46:0] twiddle4_2_366_imag;
  wire[46:0] T13654;
  wire[46:0] T13655;
  wire[46:0] T13656;
  wire[46:0] T13657;
  wire[46:0] twiddle4_2_367_imag;
  wire[46:0] T13658;
  wire[46:0] T13659;
  wire[46:0] T13660;
  wire[46:0] T13661;
  wire T13662;
  wire T13663;
  wire T13664;
  wire T13665;
  wire[46:0] T13666;
  wire[46:0] T13667;
  wire[46:0] T13668;
  wire[46:0] T13669;
  wire[46:0] twiddle4_2_368_imag;
  wire[46:0] T13670;
  wire[46:0] T13671;
  wire[46:0] T13672;
  wire[46:0] T13673;
  wire[46:0] twiddle4_2_369_imag;
  wire[46:0] T13674;
  wire[46:0] T13675;
  wire[46:0] T13676;
  wire[46:0] T13677;
  wire T13678;
  wire[46:0] T13679;
  wire[46:0] twiddle4_2_370_imag;
  wire[46:0] T13680;
  wire[46:0] T13681;
  wire[46:0] T13682;
  wire[46:0] T13683;
  wire[46:0] twiddle4_2_371_imag;
  wire[46:0] T13684;
  wire[46:0] T13685;
  wire[46:0] T13686;
  wire[46:0] T13687;
  wire T13688;
  wire T13689;
  wire[46:0] T13690;
  wire[46:0] T13691;
  wire[46:0] twiddle4_2_372_imag;
  wire[46:0] T13692;
  wire[46:0] T13693;
  wire[46:0] T13694;
  wire[46:0] T13695;
  wire[46:0] twiddle4_2_373_imag;
  wire[46:0] T13696;
  wire[46:0] T13697;
  wire[46:0] T13698;
  wire[46:0] T13699;
  wire T13700;
  wire[46:0] T13701;
  wire[46:0] twiddle4_2_374_imag;
  wire[46:0] T13702;
  wire[46:0] T13703;
  wire[46:0] T13704;
  wire[46:0] T13705;
  wire[46:0] twiddle4_2_375_imag;
  wire[46:0] T13706;
  wire[46:0] T13707;
  wire[46:0] T13708;
  wire[46:0] T13709;
  wire T13710;
  wire T13711;
  wire T13712;
  wire[46:0] T13713;
  wire[46:0] T13714;
  wire[46:0] T13715;
  wire[46:0] twiddle4_2_376_imag;
  wire[46:0] T13716;
  wire[46:0] T13717;
  wire[46:0] T13718;
  wire[46:0] T13719;
  wire[46:0] twiddle4_2_377_imag;
  wire[46:0] T13720;
  wire[46:0] T13721;
  wire[46:0] T13722;
  wire[46:0] T13723;
  wire T13724;
  wire[46:0] T13725;
  wire[46:0] twiddle4_2_378_imag;
  wire[46:0] T13726;
  wire[46:0] T13727;
  wire[46:0] T13728;
  wire[46:0] T13729;
  wire[46:0] twiddle4_2_379_imag;
  wire[46:0] T13730;
  wire[46:0] T13731;
  wire[46:0] T13732;
  wire[46:0] T13733;
  wire T13734;
  wire T13735;
  wire[46:0] T13736;
  wire[46:0] T13737;
  wire[46:0] twiddle4_2_380_imag;
  wire[46:0] T13738;
  wire[46:0] T13739;
  wire[46:0] T13740;
  wire[46:0] T13741;
  wire[46:0] twiddle4_2_381_imag;
  wire[46:0] T13742;
  wire[46:0] T13743;
  wire[46:0] T13744;
  wire[46:0] T13745;
  wire T13746;
  wire[46:0] T13747;
  wire[46:0] twiddle4_2_382_imag;
  wire[46:0] T13748;
  wire[46:0] T13749;
  wire[46:0] T13750;
  wire[46:0] T13751;
  wire[46:0] twiddle4_2_383_imag;
  wire[46:0] T13752;
  wire[46:0] T13753;
  wire[46:0] T13754;
  wire[46:0] T13755;
  wire T13756;
  wire T13757;
  wire T13758;
  wire T13759;
  wire T13760;
  wire T13761;
  wire T13762;
  wire T13763;
  wire[47:0] T13764;
  wire[46:0] T13765;
  wire[46:0] T13766;
  wire[46:0] T13767;
  wire[46:0] T13768;
  wire[46:0] T13769;
  wire[46:0] T13770;
  wire[46:0] T13771;
  wire[46:0] twiddle4_2_384_imag;
  wire[46:0] T13772;
  wire[46:0] T13773;
  wire[46:0] T13774;
  wire[46:0] T13775;
  wire[46:0] twiddle4_2_385_imag;
  wire[46:0] T13776;
  wire[46:0] T13777;
  wire[46:0] T13778;
  wire[46:0] T13779;
  wire T13780;
  wire[46:0] T13781;
  wire[46:0] twiddle4_2_386_imag;
  wire[46:0] T13782;
  wire[46:0] T13783;
  wire[46:0] T13784;
  wire[46:0] T13785;
  wire[46:0] twiddle4_2_387_imag;
  wire[46:0] T13786;
  wire[46:0] T13787;
  wire[46:0] T13788;
  wire[46:0] T13789;
  wire T13790;
  wire T13791;
  wire[46:0] T13792;
  wire[46:0] T13793;
  wire[46:0] twiddle4_2_388_imag;
  wire[46:0] T13794;
  wire[46:0] T13795;
  wire[46:0] T13796;
  wire[46:0] T13797;
  wire[46:0] twiddle4_2_389_imag;
  wire[46:0] T13798;
  wire[46:0] T13799;
  wire[46:0] T13800;
  wire[46:0] T13801;
  wire T13802;
  wire[46:0] T13803;
  wire[46:0] twiddle4_2_390_imag;
  wire[46:0] T13804;
  wire[46:0] T13805;
  wire[46:0] T13806;
  wire[46:0] T13807;
  wire[46:0] twiddle4_2_391_imag;
  wire[46:0] T13808;
  wire[46:0] T13809;
  wire[46:0] T13810;
  wire[46:0] T13811;
  wire T13812;
  wire T13813;
  wire T13814;
  wire[46:0] T13815;
  wire[46:0] T13816;
  wire[46:0] T13817;
  wire[46:0] twiddle4_2_392_imag;
  wire[46:0] T13818;
  wire[46:0] T13819;
  wire[46:0] T13820;
  wire[46:0] T13821;
  wire[46:0] twiddle4_2_393_imag;
  wire[46:0] T13822;
  wire[46:0] T13823;
  wire[46:0] T13824;
  wire[46:0] T13825;
  wire T13826;
  wire[46:0] T13827;
  wire[46:0] twiddle4_2_394_imag;
  wire[46:0] T13828;
  wire[46:0] T13829;
  wire[46:0] T13830;
  wire[46:0] T13831;
  wire[46:0] twiddle4_2_395_imag;
  wire[46:0] T13832;
  wire[46:0] T13833;
  wire[46:0] T13834;
  wire[46:0] T13835;
  wire T13836;
  wire T13837;
  wire[46:0] T13838;
  wire[46:0] T13839;
  wire[46:0] twiddle4_2_396_imag;
  wire[46:0] T13840;
  wire[46:0] T13841;
  wire[46:0] T13842;
  wire[46:0] T13843;
  wire[46:0] twiddle4_2_397_imag;
  wire[46:0] T13844;
  wire[46:0] T13845;
  wire[46:0] T13846;
  wire[46:0] T13847;
  wire T13848;
  wire[46:0] T13849;
  wire[46:0] twiddle4_2_398_imag;
  wire[46:0] T13850;
  wire[46:0] T13851;
  wire[46:0] T13852;
  wire[46:0] T13853;
  wire[46:0] twiddle4_2_399_imag;
  wire[46:0] T13854;
  wire[46:0] T13855;
  wire[46:0] T13856;
  wire[46:0] T13857;
  wire T13858;
  wire T13859;
  wire T13860;
  wire T13861;
  wire[46:0] T13862;
  wire[46:0] T13863;
  wire[46:0] T13864;
  wire[46:0] T13865;
  wire[46:0] twiddle4_2_400_imag;
  wire[46:0] T13866;
  wire[46:0] T13867;
  wire[46:0] T13868;
  wire[46:0] T13869;
  wire[46:0] twiddle4_2_401_imag;
  wire[46:0] T13870;
  wire[46:0] T13871;
  wire[46:0] T13872;
  wire[46:0] T13873;
  wire T13874;
  wire[46:0] T13875;
  wire[46:0] twiddle4_2_402_imag;
  wire[46:0] T13876;
  wire[46:0] T13877;
  wire[46:0] T13878;
  wire[46:0] T13879;
  wire[46:0] twiddle4_2_403_imag;
  wire[46:0] T13880;
  wire[46:0] T13881;
  wire[46:0] T13882;
  wire[46:0] T13883;
  wire T13884;
  wire T13885;
  wire[46:0] T13886;
  wire[46:0] T13887;
  wire[46:0] twiddle4_2_404_imag;
  wire[46:0] T13888;
  wire[46:0] T13889;
  wire[46:0] T13890;
  wire[46:0] T13891;
  wire[46:0] twiddle4_2_405_imag;
  wire[46:0] T13892;
  wire[46:0] T13893;
  wire[46:0] T13894;
  wire[46:0] T13895;
  wire T13896;
  wire[46:0] T13897;
  wire[46:0] twiddle4_2_406_imag;
  wire[46:0] T13898;
  wire[46:0] T13899;
  wire[46:0] T13900;
  wire[46:0] T13901;
  wire[46:0] twiddle4_2_407_imag;
  wire[46:0] T13902;
  wire[46:0] T13903;
  wire[46:0] T13904;
  wire[46:0] T13905;
  wire T13906;
  wire T13907;
  wire T13908;
  wire[46:0] T13909;
  wire[46:0] T13910;
  wire[46:0] T13911;
  wire[46:0] twiddle4_2_408_imag;
  wire[46:0] T13912;
  wire[46:0] T13913;
  wire[46:0] T13914;
  wire[46:0] T13915;
  wire[46:0] twiddle4_2_409_imag;
  wire[46:0] T13916;
  wire[46:0] T13917;
  wire[46:0] T13918;
  wire[46:0] T13919;
  wire T13920;
  wire[46:0] T13921;
  wire[46:0] twiddle4_2_410_imag;
  wire[46:0] T13922;
  wire[46:0] T13923;
  wire[46:0] T13924;
  wire[46:0] T13925;
  wire[46:0] twiddle4_2_411_imag;
  wire[46:0] T13926;
  wire[46:0] T13927;
  wire[46:0] T13928;
  wire[46:0] T13929;
  wire T13930;
  wire T13931;
  wire[46:0] T13932;
  wire[46:0] T13933;
  wire[46:0] twiddle4_2_412_imag;
  wire[46:0] T13934;
  wire[46:0] T13935;
  wire[46:0] T13936;
  wire[46:0] T13937;
  wire[46:0] twiddle4_2_413_imag;
  wire[46:0] T13938;
  wire[46:0] T13939;
  wire[46:0] T13940;
  wire[46:0] T13941;
  wire T13942;
  wire[46:0] T13943;
  wire[46:0] twiddle4_2_414_imag;
  wire[46:0] T13944;
  wire[46:0] T13945;
  wire[46:0] T13946;
  wire[46:0] T13947;
  wire[46:0] twiddle4_2_415_imag;
  wire[46:0] T13948;
  wire[46:0] T13949;
  wire[46:0] T13950;
  wire[46:0] T13951;
  wire T13952;
  wire T13953;
  wire T13954;
  wire T13955;
  wire T13956;
  wire[46:0] T13957;
  wire[46:0] T13958;
  wire[46:0] T13959;
  wire[46:0] T13960;
  wire[46:0] T13961;
  wire[46:0] twiddle4_2_416_imag;
  wire[46:0] T13962;
  wire[46:0] T13963;
  wire[46:0] T13964;
  wire[46:0] T13965;
  wire[46:0] twiddle4_2_417_imag;
  wire[46:0] T13966;
  wire[46:0] T13967;
  wire[46:0] T13968;
  wire[46:0] T13969;
  wire T13970;
  wire[46:0] T13971;
  wire[46:0] twiddle4_2_418_imag;
  wire[46:0] T13972;
  wire[46:0] T13973;
  wire[46:0] T13974;
  wire[46:0] T13975;
  wire[46:0] twiddle4_2_419_imag;
  wire[46:0] T13976;
  wire[46:0] T13977;
  wire[46:0] T13978;
  wire[46:0] T13979;
  wire T13980;
  wire T13981;
  wire[46:0] T13982;
  wire[46:0] T13983;
  wire[46:0] twiddle4_2_420_imag;
  wire[46:0] T13984;
  wire[46:0] T13985;
  wire[46:0] T13986;
  wire[46:0] T13987;
  wire[46:0] twiddle4_2_421_imag;
  wire[46:0] T13988;
  wire[46:0] T13989;
  wire[46:0] T13990;
  wire[46:0] T13991;
  wire T13992;
  wire[46:0] T13993;
  wire[46:0] twiddle4_2_422_imag;
  wire[46:0] T13994;
  wire[46:0] T13995;
  wire[46:0] T13996;
  wire[46:0] T13997;
  wire[46:0] twiddle4_2_423_imag;
  wire[46:0] T13998;
  wire[46:0] T13999;
  wire[46:0] T14000;
  wire[46:0] T14001;
  wire T14002;
  wire T14003;
  wire T14004;
  wire[46:0] T14005;
  wire[46:0] T14006;
  wire[46:0] T14007;
  wire[46:0] twiddle4_2_424_imag;
  wire[46:0] T14008;
  wire[46:0] T14009;
  wire[46:0] T14010;
  wire[46:0] T14011;
  wire[46:0] twiddle4_2_425_imag;
  wire[46:0] T14012;
  wire[46:0] T14013;
  wire[46:0] T14014;
  wire[46:0] T14015;
  wire T14016;
  wire[46:0] T14017;
  wire[46:0] twiddle4_2_426_imag;
  wire[46:0] T14018;
  wire[46:0] T14019;
  wire[46:0] T14020;
  wire[46:0] T14021;
  wire[46:0] twiddle4_2_427_imag;
  wire[46:0] T14022;
  wire[45:0] T14023;
  wire[45:0] T14024;
  wire T14025;
  wire[46:0] T14026;
  wire[46:0] T14027;
  wire T14028;
  wire T14029;
  wire[46:0] T14030;
  wire[46:0] T14031;
  wire[46:0] twiddle4_2_428_imag;
  wire[46:0] T14032;
  wire[45:0] T14033;
  wire[45:0] T14034;
  wire T14035;
  wire[46:0] T14036;
  wire[46:0] T14037;
  wire[46:0] twiddle4_2_429_imag;
  wire[46:0] T14038;
  wire[45:0] T14039;
  wire[45:0] T14040;
  wire T14041;
  wire[46:0] T14042;
  wire[46:0] T14043;
  wire T14044;
  wire[46:0] T14045;
  wire[46:0] twiddle4_2_430_imag;
  wire[46:0] T14046;
  wire[45:0] T14047;
  wire[45:0] T14048;
  wire T14049;
  wire[46:0] T14050;
  wire[46:0] T14051;
  wire[46:0] twiddle4_2_431_imag;
  wire[46:0] T14052;
  wire[45:0] T14053;
  wire[45:0] T14054;
  wire T14055;
  wire[46:0] T14056;
  wire[46:0] T14057;
  wire T14058;
  wire T14059;
  wire T14060;
  wire T14061;
  wire[46:0] T14062;
  wire[46:0] T14063;
  wire[46:0] T14064;
  wire[46:0] T14065;
  wire[46:0] twiddle4_2_432_imag;
  wire[46:0] T14066;
  wire[45:0] T14067;
  wire[45:0] T14068;
  wire T14069;
  wire[46:0] T14070;
  wire[46:0] T14071;
  wire[46:0] twiddle4_2_433_imag;
  wire[46:0] T14072;
  wire[45:0] T14073;
  wire[45:0] T14074;
  wire T14075;
  wire[46:0] T14076;
  wire[46:0] T14077;
  wire T14078;
  wire[46:0] T14079;
  wire[46:0] twiddle4_2_434_imag;
  wire[46:0] T14080;
  wire[45:0] T14081;
  wire[45:0] T14082;
  wire T14083;
  wire[46:0] T14084;
  wire[46:0] T14085;
  wire[46:0] twiddle4_2_435_imag;
  wire[46:0] T14086;
  wire[45:0] T14087;
  wire[45:0] T14088;
  wire T14089;
  wire[46:0] T14090;
  wire[46:0] T14091;
  wire T14092;
  wire T14093;
  wire[46:0] T14094;
  wire[46:0] T14095;
  wire[46:0] twiddle4_2_436_imag;
  wire[46:0] T14096;
  wire[45:0] T14097;
  wire[45:0] T14098;
  wire T14099;
  wire[46:0] T14100;
  wire[46:0] T14101;
  wire[46:0] twiddle4_2_437_imag;
  wire[46:0] T14102;
  wire[45:0] T14103;
  wire[45:0] T14104;
  wire T14105;
  wire[46:0] T14106;
  wire[46:0] T14107;
  wire T14108;
  wire[46:0] T14109;
  wire[46:0] twiddle4_2_438_imag;
  wire[46:0] T14110;
  wire[45:0] T14111;
  wire[45:0] T14112;
  wire T14113;
  wire[46:0] T14114;
  wire[46:0] T14115;
  wire[46:0] twiddle4_2_439_imag;
  wire[46:0] T14116;
  wire[45:0] T14117;
  wire[45:0] T14118;
  wire T14119;
  wire[46:0] T14120;
  wire[46:0] T14121;
  wire T14122;
  wire T14123;
  wire T14124;
  wire[46:0] T14125;
  wire[46:0] T14126;
  wire[46:0] T14127;
  wire[46:0] twiddle4_2_440_imag;
  wire[46:0] T14128;
  wire[45:0] T14129;
  wire[45:0] T14130;
  wire T14131;
  wire[46:0] T14132;
  wire[46:0] T14133;
  wire[46:0] twiddle4_2_441_imag;
  wire[46:0] T14134;
  wire[45:0] T14135;
  wire[45:0] T14136;
  wire T14137;
  wire[46:0] T14138;
  wire[46:0] T14139;
  wire T14140;
  wire[46:0] T14141;
  wire[46:0] twiddle4_2_442_imag;
  wire[46:0] T14142;
  wire[45:0] T14143;
  wire[45:0] T14144;
  wire T14145;
  wire[46:0] T14146;
  wire[46:0] T14147;
  wire[46:0] twiddle4_2_443_imag;
  wire[46:0] T14148;
  wire[45:0] T14149;
  wire[45:0] T14150;
  wire T14151;
  wire[46:0] T14152;
  wire[46:0] T14153;
  wire T14154;
  wire T14155;
  wire[46:0] T14156;
  wire[46:0] T14157;
  wire[46:0] twiddle4_2_444_imag;
  wire[46:0] T14158;
  wire[45:0] T14159;
  wire[45:0] T14160;
  wire T14161;
  wire[46:0] T14162;
  wire[46:0] T14163;
  wire[46:0] twiddle4_2_445_imag;
  wire[46:0] T14164;
  wire[45:0] T14165;
  wire[45:0] T14166;
  wire T14167;
  wire[46:0] T14168;
  wire[46:0] T14169;
  wire T14170;
  wire[46:0] T14171;
  wire[46:0] twiddle4_2_446_imag;
  wire[46:0] T14172;
  wire[45:0] T14173;
  wire[45:0] T14174;
  wire T14175;
  wire[46:0] T14176;
  wire[46:0] T14177;
  wire[46:0] twiddle4_2_447_imag;
  wire[46:0] T14178;
  wire[45:0] T14179;
  wire[45:0] T14180;
  wire T14181;
  wire[46:0] T14182;
  wire[46:0] T14183;
  wire T14184;
  wire T14185;
  wire T14186;
  wire T14187;
  wire T14188;
  wire T14189;
  wire[46:0] T14190;
  wire[46:0] T14191;
  wire[46:0] T14192;
  wire[46:0] T14193;
  wire[46:0] T14194;
  wire[46:0] T14195;
  wire[46:0] twiddle4_2_448_imag;
  wire[46:0] T14196;
  wire[45:0] T14197;
  wire[45:0] T14198;
  wire T14199;
  wire[46:0] T14200;
  wire[46:0] T14201;
  wire[46:0] twiddle4_2_449_imag;
  wire[46:0] T14202;
  wire[45:0] T14203;
  wire[45:0] T14204;
  wire T14205;
  wire[46:0] T14206;
  wire[46:0] T14207;
  wire T14208;
  wire[46:0] T14209;
  wire[46:0] twiddle4_2_450_imag;
  wire[46:0] T14210;
  wire[45:0] T14211;
  wire[45:0] T14212;
  wire T14213;
  wire[46:0] T14214;
  wire[46:0] T14215;
  wire[46:0] twiddle4_2_451_imag;
  wire[46:0] T14216;
  wire[45:0] T14217;
  wire[45:0] T14218;
  wire T14219;
  wire[46:0] T14220;
  wire[46:0] T14221;
  wire T14222;
  wire T14223;
  wire[46:0] T14224;
  wire[46:0] T14225;
  wire[46:0] twiddle4_2_452_imag;
  wire[46:0] T14226;
  wire[45:0] T14227;
  wire[45:0] T14228;
  wire T14229;
  wire[46:0] T14230;
  wire[46:0] T14231;
  wire[46:0] twiddle4_2_453_imag;
  wire[46:0] T14232;
  wire[45:0] T14233;
  wire[45:0] T14234;
  wire T14235;
  wire[46:0] T14236;
  wire[46:0] T14237;
  wire T14238;
  wire[46:0] T14239;
  wire[46:0] twiddle4_2_454_imag;
  wire[46:0] T14240;
  wire[45:0] T14241;
  wire[45:0] T14242;
  wire T14243;
  wire[46:0] T14244;
  wire[46:0] T14245;
  wire[46:0] twiddle4_2_455_imag;
  wire[46:0] T14246;
  wire[45:0] T14247;
  wire[45:0] T14248;
  wire T14249;
  wire[46:0] T14250;
  wire[46:0] T14251;
  wire T14252;
  wire T14253;
  wire T14254;
  wire[46:0] T14255;
  wire[46:0] T14256;
  wire[46:0] T14257;
  wire[46:0] twiddle4_2_456_imag;
  wire[46:0] T14258;
  wire[45:0] T14259;
  wire[45:0] T14260;
  wire T14261;
  wire[46:0] T14262;
  wire[46:0] T14263;
  wire[46:0] twiddle4_2_457_imag;
  wire[46:0] T14264;
  wire[45:0] T14265;
  wire[45:0] T14266;
  wire T14267;
  wire[46:0] T14268;
  wire[46:0] T14269;
  wire T14270;
  wire[46:0] T14271;
  wire[46:0] twiddle4_2_458_imag;
  wire[46:0] T14272;
  wire[45:0] T14273;
  wire[45:0] T14274;
  wire T14275;
  wire[46:0] T14276;
  wire[46:0] T14277;
  wire[46:0] twiddle4_2_459_imag;
  wire[46:0] T14278;
  wire[45:0] T14279;
  wire[45:0] T14280;
  wire T14281;
  wire[46:0] T14282;
  wire[46:0] T14283;
  wire T14284;
  wire T14285;
  wire[46:0] T14286;
  wire[46:0] T14287;
  wire[46:0] twiddle4_2_460_imag;
  wire[46:0] T14288;
  wire[45:0] T14289;
  wire[45:0] T14290;
  wire T14291;
  wire[46:0] T14292;
  wire[46:0] T14293;
  wire[46:0] twiddle4_2_461_imag;
  wire[46:0] T14294;
  wire[45:0] T14295;
  wire[45:0] T14296;
  wire T14297;
  wire[46:0] T14298;
  wire[46:0] T14299;
  wire T14300;
  wire[46:0] T14301;
  wire[46:0] twiddle4_2_462_imag;
  wire[46:0] T14302;
  wire[45:0] T14303;
  wire[45:0] T14304;
  wire T14305;
  wire[46:0] T14306;
  wire[46:0] T14307;
  wire[46:0] twiddle4_2_463_imag;
  wire[46:0] T14308;
  wire[45:0] T14309;
  wire[45:0] T14310;
  wire T14311;
  wire[46:0] T14312;
  wire[46:0] T14313;
  wire T14314;
  wire T14315;
  wire T14316;
  wire T14317;
  wire[46:0] T14318;
  wire[46:0] T14319;
  wire[46:0] T14320;
  wire[46:0] T14321;
  wire[46:0] twiddle4_2_464_imag;
  wire[46:0] T14322;
  wire[45:0] T14323;
  wire[45:0] T14324;
  wire T14325;
  wire[46:0] T14326;
  wire[46:0] T14327;
  wire[46:0] twiddle4_2_465_imag;
  wire[46:0] T14328;
  wire[45:0] T14329;
  wire[45:0] T14330;
  wire T14331;
  wire[46:0] T14332;
  wire[46:0] T14333;
  wire T14334;
  wire[46:0] T14335;
  wire[46:0] twiddle4_2_466_imag;
  wire[46:0] T14336;
  wire[45:0] T14337;
  wire[45:0] T14338;
  wire T14339;
  wire[46:0] T14340;
  wire[46:0] T14341;
  wire[46:0] twiddle4_2_467_imag;
  wire[46:0] T14342;
  wire[45:0] T14343;
  wire[45:0] T14344;
  wire T14345;
  wire[46:0] T14346;
  wire[46:0] T14347;
  wire T14348;
  wire T14349;
  wire[46:0] T14350;
  wire[46:0] T14351;
  wire[46:0] twiddle4_2_468_imag;
  wire[46:0] T14352;
  wire[45:0] T14353;
  wire[45:0] T14354;
  wire T14355;
  wire[46:0] T14356;
  wire[46:0] T14357;
  wire[46:0] twiddle4_2_469_imag;
  wire[46:0] T14358;
  wire[45:0] T14359;
  wire[45:0] T14360;
  wire T14361;
  wire[46:0] T14362;
  wire[46:0] T14363;
  wire T14364;
  wire[46:0] T14365;
  wire[46:0] twiddle4_2_470_imag;
  wire[46:0] T14366;
  wire[45:0] T14367;
  wire[45:0] T14368;
  wire T14369;
  wire[46:0] T14370;
  wire[46:0] T14371;
  wire[46:0] twiddle4_2_471_imag;
  wire[46:0] T14372;
  wire[44:0] T14373;
  wire[44:0] T14374;
  wire[1:0] T14375;
  wire T14376;
  wire[46:0] T14377;
  wire[46:0] T14378;
  wire T14379;
  wire T14380;
  wire T14381;
  wire[46:0] T14382;
  wire[46:0] T14383;
  wire[46:0] T14384;
  wire[46:0] twiddle4_2_472_imag;
  wire[46:0] T14385;
  wire[44:0] T14386;
  wire[44:0] T14387;
  wire[1:0] T14388;
  wire T14389;
  wire[46:0] T14390;
  wire[46:0] T14391;
  wire[46:0] twiddle4_2_473_imag;
  wire[46:0] T14392;
  wire[44:0] T14393;
  wire[44:0] T14394;
  wire[1:0] T14395;
  wire T14396;
  wire[46:0] T14397;
  wire[46:0] T14398;
  wire T14399;
  wire[46:0] T14400;
  wire[46:0] twiddle4_2_474_imag;
  wire[46:0] T14401;
  wire[44:0] T14402;
  wire[44:0] T14403;
  wire[1:0] T14404;
  wire T14405;
  wire[46:0] T14406;
  wire[46:0] T14407;
  wire[46:0] twiddle4_2_475_imag;
  wire[46:0] T14408;
  wire[44:0] T14409;
  wire[44:0] T14410;
  wire[1:0] T14411;
  wire T14412;
  wire[46:0] T14413;
  wire[46:0] T14414;
  wire T14415;
  wire T14416;
  wire[46:0] T14417;
  wire[46:0] T14418;
  wire[46:0] twiddle4_2_476_imag;
  wire[46:0] T14419;
  wire[44:0] T14420;
  wire[44:0] T14421;
  wire[1:0] T14422;
  wire T14423;
  wire[46:0] T14424;
  wire[46:0] T14425;
  wire[46:0] twiddle4_2_477_imag;
  wire[46:0] T14426;
  wire[44:0] T14427;
  wire[44:0] T14428;
  wire[1:0] T14429;
  wire T14430;
  wire[46:0] T14431;
  wire[46:0] T14432;
  wire T14433;
  wire[46:0] T14434;
  wire[46:0] twiddle4_2_478_imag;
  wire[46:0] T14435;
  wire[44:0] T14436;
  wire[44:0] T14437;
  wire[1:0] T14438;
  wire T14439;
  wire[46:0] T14440;
  wire[46:0] T14441;
  wire[46:0] twiddle4_2_479_imag;
  wire[46:0] T14442;
  wire[44:0] T14443;
  wire[44:0] T14444;
  wire[1:0] T14445;
  wire T14446;
  wire[46:0] T14447;
  wire[46:0] T14448;
  wire T14449;
  wire T14450;
  wire T14451;
  wire T14452;
  wire T14453;
  wire[46:0] T14454;
  wire[46:0] T14455;
  wire[46:0] T14456;
  wire[46:0] T14457;
  wire[46:0] T14458;
  wire[46:0] twiddle4_2_480_imag;
  wire[46:0] T14459;
  wire[44:0] T14460;
  wire[44:0] T14461;
  wire[1:0] T14462;
  wire T14463;
  wire[46:0] T14464;
  wire[46:0] T14465;
  wire[46:0] twiddle4_2_481_imag;
  wire[46:0] T14466;
  wire[44:0] T14467;
  wire[44:0] T14468;
  wire[1:0] T14469;
  wire T14470;
  wire[46:0] T14471;
  wire[46:0] T14472;
  wire T14473;
  wire[46:0] T14474;
  wire[46:0] twiddle4_2_482_imag;
  wire[46:0] T14475;
  wire[44:0] T14476;
  wire[44:0] T14477;
  wire[1:0] T14478;
  wire T14479;
  wire[46:0] T14480;
  wire[46:0] T14481;
  wire[46:0] twiddle4_2_483_imag;
  wire[46:0] T14482;
  wire[44:0] T14483;
  wire[44:0] T14484;
  wire[1:0] T14485;
  wire T14486;
  wire[46:0] T14487;
  wire[46:0] T14488;
  wire T14489;
  wire T14490;
  wire[46:0] T14491;
  wire[46:0] T14492;
  wire[46:0] twiddle4_2_484_imag;
  wire[46:0] T14493;
  wire[44:0] T14494;
  wire[44:0] T14495;
  wire[1:0] T14496;
  wire T14497;
  wire[46:0] T14498;
  wire[46:0] T14499;
  wire[46:0] twiddle4_2_485_imag;
  wire[46:0] T14500;
  wire[44:0] T14501;
  wire[44:0] T14502;
  wire[1:0] T14503;
  wire T14504;
  wire[46:0] T14505;
  wire[46:0] T14506;
  wire T14507;
  wire[46:0] T14508;
  wire[46:0] twiddle4_2_486_imag;
  wire[46:0] T14509;
  wire[44:0] T14510;
  wire[44:0] T14511;
  wire[1:0] T14512;
  wire T14513;
  wire[46:0] T14514;
  wire[46:0] T14515;
  wire[46:0] twiddle4_2_487_imag;
  wire[46:0] T14516;
  wire[44:0] T14517;
  wire[44:0] T14518;
  wire[1:0] T14519;
  wire T14520;
  wire[46:0] T14521;
  wire[46:0] T14522;
  wire T14523;
  wire T14524;
  wire T14525;
  wire[46:0] T14526;
  wire[46:0] T14527;
  wire[46:0] T14528;
  wire[46:0] twiddle4_2_488_imag;
  wire[46:0] T14529;
  wire[44:0] T14530;
  wire[44:0] T14531;
  wire[1:0] T14532;
  wire T14533;
  wire[46:0] T14534;
  wire[46:0] T14535;
  wire[46:0] twiddle4_2_489_imag;
  wire[46:0] T14536;
  wire[44:0] T14537;
  wire[44:0] T14538;
  wire[1:0] T14539;
  wire T14540;
  wire[46:0] T14541;
  wire[46:0] T14542;
  wire T14543;
  wire[46:0] T14544;
  wire[46:0] twiddle4_2_490_imag;
  wire[46:0] T14545;
  wire[44:0] T14546;
  wire[44:0] T14547;
  wire[1:0] T14548;
  wire T14549;
  wire[46:0] T14550;
  wire[46:0] T14551;
  wire[46:0] twiddle4_2_491_imag;
  wire[46:0] T14552;
  wire[44:0] T14553;
  wire[44:0] T14554;
  wire[1:0] T14555;
  wire T14556;
  wire[46:0] T14557;
  wire[46:0] T14558;
  wire T14559;
  wire T14560;
  wire[46:0] T14561;
  wire[46:0] T14562;
  wire[46:0] twiddle4_2_492_imag;
  wire[46:0] T14563;
  wire[43:0] T14564;
  wire[43:0] T14565;
  wire[2:0] T14566;
  wire T14567;
  wire[46:0] T14568;
  wire[46:0] T14569;
  wire[46:0] twiddle4_2_493_imag;
  wire[46:0] T14570;
  wire[43:0] T14571;
  wire[43:0] T14572;
  wire[2:0] T14573;
  wire T14574;
  wire[46:0] T14575;
  wire[46:0] T14576;
  wire T14577;
  wire[46:0] T14578;
  wire[46:0] twiddle4_2_494_imag;
  wire[46:0] T14579;
  wire[43:0] T14580;
  wire[43:0] T14581;
  wire[2:0] T14582;
  wire T14583;
  wire[46:0] T14584;
  wire[46:0] T14585;
  wire[46:0] twiddle4_2_495_imag;
  wire[46:0] T14586;
  wire[43:0] T14587;
  wire[43:0] T14588;
  wire[2:0] T14589;
  wire T14590;
  wire[46:0] T14591;
  wire[46:0] T14592;
  wire T14593;
  wire T14594;
  wire T14595;
  wire T14596;
  wire[46:0] T14597;
  wire[46:0] T14598;
  wire[46:0] T14599;
  wire[46:0] T14600;
  wire[46:0] twiddle4_2_496_imag;
  wire[46:0] T14601;
  wire[43:0] T14602;
  wire[43:0] T14603;
  wire[2:0] T14604;
  wire T14605;
  wire[46:0] T14606;
  wire[46:0] T14607;
  wire[46:0] twiddle4_2_497_imag;
  wire[46:0] T14608;
  wire[43:0] T14609;
  wire[43:0] T14610;
  wire[2:0] T14611;
  wire T14612;
  wire[46:0] T14613;
  wire[46:0] T14614;
  wire T14615;
  wire[46:0] T14616;
  wire[46:0] twiddle4_2_498_imag;
  wire[46:0] T14617;
  wire[43:0] T14618;
  wire[43:0] T14619;
  wire[2:0] T14620;
  wire T14621;
  wire[46:0] T14622;
  wire[46:0] T14623;
  wire[46:0] twiddle4_2_499_imag;
  wire[46:0] T14624;
  wire[43:0] T14625;
  wire[43:0] T14626;
  wire[2:0] T14627;
  wire T14628;
  wire[46:0] T14629;
  wire[46:0] T14630;
  wire T14631;
  wire T14632;
  wire[46:0] T14633;
  wire[46:0] T14634;
  wire[46:0] twiddle4_2_500_imag;
  wire[46:0] T14635;
  wire[43:0] T14636;
  wire[43:0] T14637;
  wire[2:0] T14638;
  wire T14639;
  wire[46:0] T14640;
  wire[46:0] T14641;
  wire[46:0] twiddle4_2_501_imag;
  wire[46:0] T14642;
  wire[43:0] T14643;
  wire[43:0] T14644;
  wire[2:0] T14645;
  wire T14646;
  wire[46:0] T14647;
  wire[46:0] T14648;
  wire T14649;
  wire[46:0] T14650;
  wire[46:0] twiddle4_2_502_imag;
  wire[46:0] T14651;
  wire[42:0] T14652;
  wire[42:0] T14653;
  wire[3:0] T14654;
  wire T14655;
  wire[46:0] T14656;
  wire[46:0] T14657;
  wire[46:0] twiddle4_2_503_imag;
  wire[46:0] T14658;
  wire[42:0] T14659;
  wire[42:0] T14660;
  wire[3:0] T14661;
  wire T14662;
  wire[46:0] T14663;
  wire[46:0] T14664;
  wire T14665;
  wire T14666;
  wire T14667;
  wire[46:0] T14668;
  wire[46:0] T14669;
  wire[46:0] T14670;
  wire[46:0] twiddle4_2_504_imag;
  wire[46:0] T14671;
  wire[42:0] T14672;
  wire[42:0] T14673;
  wire[3:0] T14674;
  wire T14675;
  wire[46:0] T14676;
  wire[46:0] T14677;
  wire[46:0] twiddle4_2_505_imag;
  wire[46:0] T14678;
  wire[42:0] T14679;
  wire[42:0] T14680;
  wire[3:0] T14681;
  wire T14682;
  wire[46:0] T14683;
  wire[46:0] T14684;
  wire T14685;
  wire[46:0] T14686;
  wire[46:0] twiddle4_2_506_imag;
  wire[46:0] T14687;
  wire[42:0] T14688;
  wire[42:0] T14689;
  wire[3:0] T14690;
  wire T14691;
  wire[46:0] T14692;
  wire[46:0] T14693;
  wire[46:0] twiddle4_2_507_imag;
  wire[46:0] T14694;
  wire[41:0] T14695;
  wire[41:0] T14696;
  wire[4:0] T14697;
  wire T14698;
  wire[46:0] T14699;
  wire[46:0] T14700;
  wire T14701;
  wire T14702;
  wire[46:0] T14703;
  wire[46:0] T14704;
  wire[46:0] twiddle4_2_508_imag;
  wire[46:0] T14705;
  wire[41:0] T14706;
  wire[41:0] T14707;
  wire[4:0] T14708;
  wire T14709;
  wire[46:0] T14710;
  wire[46:0] T14711;
  wire[46:0] twiddle4_2_509_imag;
  wire[46:0] T14712;
  wire[41:0] T14713;
  wire[41:0] T14714;
  wire[4:0] T14715;
  wire T14716;
  wire[46:0] T14717;
  wire[46:0] T14718;
  wire T14719;
  wire[46:0] T14720;
  wire[46:0] twiddle4_2_510_imag;
  wire[46:0] T14721;
  wire[40:0] T14722;
  wire[40:0] T14723;
  wire[5:0] T14724;
  wire T14725;
  wire[46:0] T14726;
  wire[46:0] T14727;
  wire[46:0] twiddle4_2_511_imag;
  wire[46:0] T14728;
  wire[39:0] T14729;
  wire[39:0] T14730;
  wire[6:0] T14731;
  wire T14732;
  wire[46:0] T14733;
  wire[46:0] T14734;
  wire T14735;
  wire T14736;
  wire T14737;
  wire T14738;
  wire T14739;
  wire T14740;
  wire T14741;
  wire T14742;
  wire T14743;
  wire T14744;
  wire[15:0] T14745;
  wire[47:0] T14746;
  wire[47:0] T14747;
  wire[47:0] T14748;
  wire[47:0] T14749;
  wire[47:0] T14750;
  wire[47:0] T14751;
  wire[47:0] T14752;
  wire[47:0] T14753;
  wire[47:0] T14754;
  wire[47:0] twiddle4_2_0_real;
  wire[47:0] T14755;
  wire[16:0] T14756;
  wire[16:0] T14757;
  wire[30:0] T14758;
  wire T14759;
  wire[47:0] T14760;
  wire[47:0] T14761;
  wire[47:0] T14762;
  wire[46:0] twiddle4_2_1_real;
  wire[46:0] T14763;
  wire[39:0] T14764;
  wire[39:0] T14765;
  wire[6:0] T14766;
  wire T14767;
  wire[46:0] T14768;
  wire[46:0] T14769;
  wire T14770;
  wire T14771;
  wire[47:0] T14772;
  wire[46:0] T14773;
  wire[46:0] twiddle4_2_2_real;
  wire[46:0] T14774;
  wire[40:0] T14775;
  wire[40:0] T14776;
  wire[5:0] T14777;
  wire T14778;
  wire[46:0] T14779;
  wire[46:0] T14780;
  wire[46:0] twiddle4_2_3_real;
  wire[46:0] T14781;
  wire[41:0] T14782;
  wire[41:0] T14783;
  wire[4:0] T14784;
  wire T14785;
  wire[46:0] T14786;
  wire[46:0] T14787;
  wire T14788;
  wire T14789;
  wire T14790;
  wire[47:0] T14791;
  wire[46:0] T14792;
  wire[46:0] T14793;
  wire[46:0] twiddle4_2_4_real;
  wire[46:0] T14794;
  wire[41:0] T14795;
  wire[41:0] T14796;
  wire[4:0] T14797;
  wire T14798;
  wire[46:0] T14799;
  wire[46:0] T14800;
  wire[46:0] twiddle4_2_5_real;
  wire[46:0] T14801;
  wire[41:0] T14802;
  wire[41:0] T14803;
  wire[4:0] T14804;
  wire T14805;
  wire[46:0] T14806;
  wire[46:0] T14807;
  wire T14808;
  wire[46:0] T14809;
  wire[46:0] twiddle4_2_6_real;
  wire[46:0] T14810;
  wire[42:0] T14811;
  wire[42:0] T14812;
  wire[3:0] T14813;
  wire T14814;
  wire[46:0] T14815;
  wire[46:0] T14816;
  wire[46:0] twiddle4_2_7_real;
  wire[46:0] T14817;
  wire[42:0] T14818;
  wire[42:0] T14819;
  wire[3:0] T14820;
  wire T14821;
  wire[46:0] T14822;
  wire[46:0] T14823;
  wire T14824;
  wire T14825;
  wire T14826;
  wire T14827;
  wire[47:0] T14828;
  wire[46:0] T14829;
  wire[46:0] T14830;
  wire[46:0] T14831;
  wire[46:0] twiddle4_2_8_real;
  wire[46:0] T14832;
  wire[42:0] T14833;
  wire[42:0] T14834;
  wire[3:0] T14835;
  wire T14836;
  wire[46:0] T14837;
  wire[46:0] T14838;
  wire[46:0] twiddle4_2_9_real;
  wire[46:0] T14839;
  wire[42:0] T14840;
  wire[42:0] T14841;
  wire[3:0] T14842;
  wire T14843;
  wire[46:0] T14844;
  wire[46:0] T14845;
  wire T14846;
  wire[46:0] T14847;
  wire[46:0] twiddle4_2_10_real;
  wire[46:0] T14848;
  wire[42:0] T14849;
  wire[42:0] T14850;
  wire[3:0] T14851;
  wire T14852;
  wire[46:0] T14853;
  wire[46:0] T14854;
  wire[46:0] twiddle4_2_11_real;
  wire[46:0] T14855;
  wire[43:0] T14856;
  wire[43:0] T14857;
  wire[2:0] T14858;
  wire T14859;
  wire[46:0] T14860;
  wire[46:0] T14861;
  wire T14862;
  wire T14863;
  wire[46:0] T14864;
  wire[46:0] T14865;
  wire[46:0] twiddle4_2_12_real;
  wire[46:0] T14866;
  wire[43:0] T14867;
  wire[43:0] T14868;
  wire[2:0] T14869;
  wire T14870;
  wire[46:0] T14871;
  wire[46:0] T14872;
  wire[46:0] twiddle4_2_13_real;
  wire[46:0] T14873;
  wire[43:0] T14874;
  wire[43:0] T14875;
  wire[2:0] T14876;
  wire T14877;
  wire[46:0] T14878;
  wire[46:0] T14879;
  wire T14880;
  wire[46:0] T14881;
  wire[46:0] twiddle4_2_14_real;
  wire[46:0] T14882;
  wire[43:0] T14883;
  wire[43:0] T14884;
  wire[2:0] T14885;
  wire T14886;
  wire[46:0] T14887;
  wire[46:0] T14888;
  wire[46:0] twiddle4_2_15_real;
  wire[46:0] T14889;
  wire[43:0] T14890;
  wire[43:0] T14891;
  wire[2:0] T14892;
  wire T14893;
  wire[46:0] T14894;
  wire[46:0] T14895;
  wire T14896;
  wire T14897;
  wire T14898;
  wire T14899;
  wire T14900;
  wire[47:0] T14901;
  wire[46:0] T14902;
  wire[46:0] T14903;
  wire[46:0] T14904;
  wire[46:0] T14905;
  wire[46:0] twiddle4_2_16_real;
  wire[46:0] T14906;
  wire[43:0] T14907;
  wire[43:0] T14908;
  wire[2:0] T14909;
  wire T14910;
  wire[46:0] T14911;
  wire[46:0] T14912;
  wire[46:0] twiddle4_2_17_real;
  wire[46:0] T14913;
  wire[43:0] T14914;
  wire[43:0] T14915;
  wire[2:0] T14916;
  wire T14917;
  wire[46:0] T14918;
  wire[46:0] T14919;
  wire T14920;
  wire[46:0] T14921;
  wire[46:0] twiddle4_2_18_real;
  wire[46:0] T14922;
  wire[43:0] T14923;
  wire[43:0] T14924;
  wire[2:0] T14925;
  wire T14926;
  wire[46:0] T14927;
  wire[46:0] T14928;
  wire[46:0] twiddle4_2_19_real;
  wire[46:0] T14929;
  wire[43:0] T14930;
  wire[43:0] T14931;
  wire[2:0] T14932;
  wire T14933;
  wire[46:0] T14934;
  wire[46:0] T14935;
  wire T14936;
  wire T14937;
  wire[46:0] T14938;
  wire[46:0] T14939;
  wire[46:0] twiddle4_2_20_real;
  wire[46:0] T14940;
  wire[43:0] T14941;
  wire[43:0] T14942;
  wire[2:0] T14943;
  wire T14944;
  wire[46:0] T14945;
  wire[46:0] T14946;
  wire[46:0] twiddle4_2_21_real;
  wire[46:0] T14947;
  wire[44:0] T14948;
  wire[44:0] T14949;
  wire[1:0] T14950;
  wire T14951;
  wire[46:0] T14952;
  wire[46:0] T14953;
  wire T14954;
  wire[46:0] T14955;
  wire[46:0] twiddle4_2_22_real;
  wire[46:0] T14956;
  wire[44:0] T14957;
  wire[44:0] T14958;
  wire[1:0] T14959;
  wire T14960;
  wire[46:0] T14961;
  wire[46:0] T14962;
  wire[46:0] twiddle4_2_23_real;
  wire[46:0] T14963;
  wire[44:0] T14964;
  wire[44:0] T14965;
  wire[1:0] T14966;
  wire T14967;
  wire[46:0] T14968;
  wire[46:0] T14969;
  wire T14970;
  wire T14971;
  wire T14972;
  wire[46:0] T14973;
  wire[46:0] T14974;
  wire[46:0] T14975;
  wire[46:0] twiddle4_2_24_real;
  wire[46:0] T14976;
  wire[44:0] T14977;
  wire[44:0] T14978;
  wire[1:0] T14979;
  wire T14980;
  wire[46:0] T14981;
  wire[46:0] T14982;
  wire[46:0] twiddle4_2_25_real;
  wire[46:0] T14983;
  wire[44:0] T14984;
  wire[44:0] T14985;
  wire[1:0] T14986;
  wire T14987;
  wire[46:0] T14988;
  wire[46:0] T14989;
  wire T14990;
  wire[46:0] T14991;
  wire[46:0] twiddle4_2_26_real;
  wire[46:0] T14992;
  wire[44:0] T14993;
  wire[44:0] T14994;
  wire[1:0] T14995;
  wire T14996;
  wire[46:0] T14997;
  wire[46:0] T14998;
  wire[46:0] twiddle4_2_27_real;
  wire[46:0] T14999;
  wire[44:0] T15000;
  wire[44:0] T15001;
  wire[1:0] T15002;
  wire T15003;
  wire[46:0] T15004;
  wire[46:0] T15005;
  wire T15006;
  wire T15007;
  wire[46:0] T15008;
  wire[46:0] T15009;
  wire[46:0] twiddle4_2_28_real;
  wire[46:0] T15010;
  wire[44:0] T15011;
  wire[44:0] T15012;
  wire[1:0] T15013;
  wire T15014;
  wire[46:0] T15015;
  wire[46:0] T15016;
  wire[46:0] twiddle4_2_29_real;
  wire[46:0] T15017;
  wire[44:0] T15018;
  wire[44:0] T15019;
  wire[1:0] T15020;
  wire T15021;
  wire[46:0] T15022;
  wire[46:0] T15023;
  wire T15024;
  wire[46:0] T15025;
  wire[46:0] twiddle4_2_30_real;
  wire[46:0] T15026;
  wire[44:0] T15027;
  wire[44:0] T15028;
  wire[1:0] T15029;
  wire T15030;
  wire[46:0] T15031;
  wire[46:0] T15032;
  wire[46:0] twiddle4_2_31_real;
  wire[46:0] T15033;
  wire[44:0] T15034;
  wire[44:0] T15035;
  wire[1:0] T15036;
  wire T15037;
  wire[46:0] T15038;
  wire[46:0] T15039;
  wire T15040;
  wire T15041;
  wire T15042;
  wire T15043;
  wire T15044;
  wire T15045;
  wire[47:0] T15046;
  wire[46:0] T15047;
  wire[46:0] T15048;
  wire[46:0] T15049;
  wire[46:0] T15050;
  wire[46:0] T15051;
  wire[46:0] twiddle4_2_32_real;
  wire[46:0] T15052;
  wire[44:0] T15053;
  wire[44:0] T15054;
  wire[1:0] T15055;
  wire T15056;
  wire[46:0] T15057;
  wire[46:0] T15058;
  wire[46:0] twiddle4_2_33_real;
  wire[46:0] T15059;
  wire[44:0] T15060;
  wire[44:0] T15061;
  wire[1:0] T15062;
  wire T15063;
  wire[46:0] T15064;
  wire[46:0] T15065;
  wire T15066;
  wire[46:0] T15067;
  wire[46:0] twiddle4_2_34_real;
  wire[46:0] T15068;
  wire[44:0] T15069;
  wire[44:0] T15070;
  wire[1:0] T15071;
  wire T15072;
  wire[46:0] T15073;
  wire[46:0] T15074;
  wire[46:0] twiddle4_2_35_real;
  wire[46:0] T15075;
  wire[44:0] T15076;
  wire[44:0] T15077;
  wire[1:0] T15078;
  wire T15079;
  wire[46:0] T15080;
  wire[46:0] T15081;
  wire T15082;
  wire T15083;
  wire[46:0] T15084;
  wire[46:0] T15085;
  wire[46:0] twiddle4_2_36_real;
  wire[46:0] T15086;
  wire[44:0] T15087;
  wire[44:0] T15088;
  wire[1:0] T15089;
  wire T15090;
  wire[46:0] T15091;
  wire[46:0] T15092;
  wire[46:0] twiddle4_2_37_real;
  wire[46:0] T15093;
  wire[44:0] T15094;
  wire[44:0] T15095;
  wire[1:0] T15096;
  wire T15097;
  wire[46:0] T15098;
  wire[46:0] T15099;
  wire T15100;
  wire[46:0] T15101;
  wire[46:0] twiddle4_2_38_real;
  wire[46:0] T15102;
  wire[44:0] T15103;
  wire[44:0] T15104;
  wire[1:0] T15105;
  wire T15106;
  wire[46:0] T15107;
  wire[46:0] T15108;
  wire[46:0] twiddle4_2_39_real;
  wire[46:0] T15109;
  wire[44:0] T15110;
  wire[44:0] T15111;
  wire[1:0] T15112;
  wire T15113;
  wire[46:0] T15114;
  wire[46:0] T15115;
  wire T15116;
  wire T15117;
  wire T15118;
  wire[46:0] T15119;
  wire[46:0] T15120;
  wire[46:0] T15121;
  wire[46:0] twiddle4_2_40_real;
  wire[46:0] T15122;
  wire[44:0] T15123;
  wire[44:0] T15124;
  wire[1:0] T15125;
  wire T15126;
  wire[46:0] T15127;
  wire[46:0] T15128;
  wire[46:0] twiddle4_2_41_real;
  wire[46:0] T15129;
  wire[44:0] T15130;
  wire[44:0] T15131;
  wire[1:0] T15132;
  wire T15133;
  wire[46:0] T15134;
  wire[46:0] T15135;
  wire T15136;
  wire[46:0] T15137;
  wire[46:0] twiddle4_2_42_real;
  wire[46:0] T15138;
  wire[45:0] T15139;
  wire[45:0] T15140;
  wire T15141;
  wire[46:0] T15142;
  wire[46:0] T15143;
  wire[46:0] twiddle4_2_43_real;
  wire[46:0] T15144;
  wire[45:0] T15145;
  wire[45:0] T15146;
  wire T15147;
  wire[46:0] T15148;
  wire[46:0] T15149;
  wire T15150;
  wire T15151;
  wire[46:0] T15152;
  wire[46:0] T15153;
  wire[46:0] twiddle4_2_44_real;
  wire[46:0] T15154;
  wire[45:0] T15155;
  wire[45:0] T15156;
  wire T15157;
  wire[46:0] T15158;
  wire[46:0] T15159;
  wire[46:0] twiddle4_2_45_real;
  wire[46:0] T15160;
  wire[45:0] T15161;
  wire[45:0] T15162;
  wire T15163;
  wire[46:0] T15164;
  wire[46:0] T15165;
  wire T15166;
  wire[46:0] T15167;
  wire[46:0] twiddle4_2_46_real;
  wire[46:0] T15168;
  wire[45:0] T15169;
  wire[45:0] T15170;
  wire T15171;
  wire[46:0] T15172;
  wire[46:0] T15173;
  wire[46:0] twiddle4_2_47_real;
  wire[46:0] T15174;
  wire[45:0] T15175;
  wire[45:0] T15176;
  wire T15177;
  wire[46:0] T15178;
  wire[46:0] T15179;
  wire T15180;
  wire T15181;
  wire T15182;
  wire T15183;
  wire[46:0] T15184;
  wire[46:0] T15185;
  wire[46:0] T15186;
  wire[46:0] T15187;
  wire[46:0] twiddle4_2_48_real;
  wire[46:0] T15188;
  wire[45:0] T15189;
  wire[45:0] T15190;
  wire T15191;
  wire[46:0] T15192;
  wire[46:0] T15193;
  wire[46:0] twiddle4_2_49_real;
  wire[46:0] T15194;
  wire[45:0] T15195;
  wire[45:0] T15196;
  wire T15197;
  wire[46:0] T15198;
  wire[46:0] T15199;
  wire T15200;
  wire[46:0] T15201;
  wire[46:0] twiddle4_2_50_real;
  wire[46:0] T15202;
  wire[45:0] T15203;
  wire[45:0] T15204;
  wire T15205;
  wire[46:0] T15206;
  wire[46:0] T15207;
  wire[46:0] twiddle4_2_51_real;
  wire[46:0] T15208;
  wire[45:0] T15209;
  wire[45:0] T15210;
  wire T15211;
  wire[46:0] T15212;
  wire[46:0] T15213;
  wire T15214;
  wire T15215;
  wire[46:0] T15216;
  wire[46:0] T15217;
  wire[46:0] twiddle4_2_52_real;
  wire[46:0] T15218;
  wire[45:0] T15219;
  wire[45:0] T15220;
  wire T15221;
  wire[46:0] T15222;
  wire[46:0] T15223;
  wire[46:0] twiddle4_2_53_real;
  wire[46:0] T15224;
  wire[45:0] T15225;
  wire[45:0] T15226;
  wire T15227;
  wire[46:0] T15228;
  wire[46:0] T15229;
  wire T15230;
  wire[46:0] T15231;
  wire[46:0] twiddle4_2_54_real;
  wire[46:0] T15232;
  wire[45:0] T15233;
  wire[45:0] T15234;
  wire T15235;
  wire[46:0] T15236;
  wire[46:0] T15237;
  wire[46:0] twiddle4_2_55_real;
  wire[46:0] T15238;
  wire[45:0] T15239;
  wire[45:0] T15240;
  wire T15241;
  wire[46:0] T15242;
  wire[46:0] T15243;
  wire T15244;
  wire T15245;
  wire T15246;
  wire[46:0] T15247;
  wire[46:0] T15248;
  wire[46:0] T15249;
  wire[46:0] twiddle4_2_56_real;
  wire[46:0] T15250;
  wire[45:0] T15251;
  wire[45:0] T15252;
  wire T15253;
  wire[46:0] T15254;
  wire[46:0] T15255;
  wire[46:0] twiddle4_2_57_real;
  wire[46:0] T15256;
  wire[45:0] T15257;
  wire[45:0] T15258;
  wire T15259;
  wire[46:0] T15260;
  wire[46:0] T15261;
  wire T15262;
  wire[46:0] T15263;
  wire[46:0] twiddle4_2_58_real;
  wire[46:0] T15264;
  wire[45:0] T15265;
  wire[45:0] T15266;
  wire T15267;
  wire[46:0] T15268;
  wire[46:0] T15269;
  wire[46:0] twiddle4_2_59_real;
  wire[46:0] T15270;
  wire[45:0] T15271;
  wire[45:0] T15272;
  wire T15273;
  wire[46:0] T15274;
  wire[46:0] T15275;
  wire T15276;
  wire T15277;
  wire[46:0] T15278;
  wire[46:0] T15279;
  wire[46:0] twiddle4_2_60_real;
  wire[46:0] T15280;
  wire[45:0] T15281;
  wire[45:0] T15282;
  wire T15283;
  wire[46:0] T15284;
  wire[46:0] T15285;
  wire[46:0] twiddle4_2_61_real;
  wire[46:0] T15286;
  wire[45:0] T15287;
  wire[45:0] T15288;
  wire T15289;
  wire[46:0] T15290;
  wire[46:0] T15291;
  wire T15292;
  wire[46:0] T15293;
  wire[46:0] twiddle4_2_62_real;
  wire[46:0] T15294;
  wire[45:0] T15295;
  wire[45:0] T15296;
  wire T15297;
  wire[46:0] T15298;
  wire[46:0] T15299;
  wire[46:0] twiddle4_2_63_real;
  wire[46:0] T15300;
  wire[45:0] T15301;
  wire[45:0] T15302;
  wire T15303;
  wire[46:0] T15304;
  wire[46:0] T15305;
  wire T15306;
  wire T15307;
  wire T15308;
  wire T15309;
  wire T15310;
  wire T15311;
  wire T15312;
  wire[47:0] T15313;
  wire[46:0] T15314;
  wire[46:0] T15315;
  wire[46:0] T15316;
  wire[46:0] T15317;
  wire[46:0] T15318;
  wire[46:0] T15319;
  wire[46:0] twiddle4_2_64_real;
  wire[46:0] T15320;
  wire[45:0] T15321;
  wire[45:0] T15322;
  wire T15323;
  wire[46:0] T15324;
  wire[46:0] T15325;
  wire[46:0] twiddle4_2_65_real;
  wire[46:0] T15326;
  wire[45:0] T15327;
  wire[45:0] T15328;
  wire T15329;
  wire[46:0] T15330;
  wire[46:0] T15331;
  wire T15332;
  wire[46:0] T15333;
  wire[46:0] twiddle4_2_66_real;
  wire[46:0] T15334;
  wire[45:0] T15335;
  wire[45:0] T15336;
  wire T15337;
  wire[46:0] T15338;
  wire[46:0] T15339;
  wire[46:0] twiddle4_2_67_real;
  wire[46:0] T15340;
  wire[45:0] T15341;
  wire[45:0] T15342;
  wire T15343;
  wire[46:0] T15344;
  wire[46:0] T15345;
  wire T15346;
  wire T15347;
  wire[46:0] T15348;
  wire[46:0] T15349;
  wire[46:0] twiddle4_2_68_real;
  wire[46:0] T15350;
  wire[45:0] T15351;
  wire[45:0] T15352;
  wire T15353;
  wire[46:0] T15354;
  wire[46:0] T15355;
  wire[46:0] twiddle4_2_69_real;
  wire[46:0] T15356;
  wire[45:0] T15357;
  wire[45:0] T15358;
  wire T15359;
  wire[46:0] T15360;
  wire[46:0] T15361;
  wire T15362;
  wire[46:0] T15363;
  wire[46:0] twiddle4_2_70_real;
  wire[46:0] T15364;
  wire[45:0] T15365;
  wire[45:0] T15366;
  wire T15367;
  wire[46:0] T15368;
  wire[46:0] T15369;
  wire[46:0] twiddle4_2_71_real;
  wire[46:0] T15370;
  wire[45:0] T15371;
  wire[45:0] T15372;
  wire T15373;
  wire[46:0] T15374;
  wire[46:0] T15375;
  wire T15376;
  wire T15377;
  wire T15378;
  wire[46:0] T15379;
  wire[46:0] T15380;
  wire[46:0] T15381;
  wire[46:0] twiddle4_2_72_real;
  wire[46:0] T15382;
  wire[45:0] T15383;
  wire[45:0] T15384;
  wire T15385;
  wire[46:0] T15386;
  wire[46:0] T15387;
  wire[46:0] twiddle4_2_73_real;
  wire[46:0] T15388;
  wire[45:0] T15389;
  wire[45:0] T15390;
  wire T15391;
  wire[46:0] T15392;
  wire[46:0] T15393;
  wire T15394;
  wire[46:0] T15395;
  wire[46:0] twiddle4_2_74_real;
  wire[46:0] T15396;
  wire[45:0] T15397;
  wire[45:0] T15398;
  wire T15399;
  wire[46:0] T15400;
  wire[46:0] T15401;
  wire[46:0] twiddle4_2_75_real;
  wire[46:0] T15402;
  wire[45:0] T15403;
  wire[45:0] T15404;
  wire T15405;
  wire[46:0] T15406;
  wire[46:0] T15407;
  wire T15408;
  wire T15409;
  wire[46:0] T15410;
  wire[46:0] T15411;
  wire[46:0] twiddle4_2_76_real;
  wire[46:0] T15412;
  wire[45:0] T15413;
  wire[45:0] T15414;
  wire T15415;
  wire[46:0] T15416;
  wire[46:0] T15417;
  wire[46:0] twiddle4_2_77_real;
  wire[46:0] T15418;
  wire[45:0] T15419;
  wire[45:0] T15420;
  wire T15421;
  wire[46:0] T15422;
  wire[46:0] T15423;
  wire T15424;
  wire[46:0] T15425;
  wire[46:0] twiddle4_2_78_real;
  wire[46:0] T15426;
  wire[45:0] T15427;
  wire[45:0] T15428;
  wire T15429;
  wire[46:0] T15430;
  wire[46:0] T15431;
  wire[46:0] twiddle4_2_79_real;
  wire[46:0] T15432;
  wire[45:0] T15433;
  wire[45:0] T15434;
  wire T15435;
  wire[46:0] T15436;
  wire[46:0] T15437;
  wire T15438;
  wire T15439;
  wire T15440;
  wire T15441;
  wire[46:0] T15442;
  wire[46:0] T15443;
  wire[46:0] T15444;
  wire[46:0] T15445;
  wire[46:0] twiddle4_2_80_real;
  wire[46:0] T15446;
  wire[45:0] T15447;
  wire[45:0] T15448;
  wire T15449;
  wire[46:0] T15450;
  wire[46:0] T15451;
  wire[46:0] twiddle4_2_81_real;
  wire[46:0] T15452;
  wire[45:0] T15453;
  wire[45:0] T15454;
  wire T15455;
  wire[46:0] T15456;
  wire[46:0] T15457;
  wire T15458;
  wire[46:0] T15459;
  wire[46:0] twiddle4_2_82_real;
  wire[46:0] T15460;
  wire[45:0] T15461;
  wire[45:0] T15462;
  wire T15463;
  wire[46:0] T15464;
  wire[46:0] T15465;
  wire[46:0] twiddle4_2_83_real;
  wire[46:0] T15466;
  wire[45:0] T15467;
  wire[45:0] T15468;
  wire T15469;
  wire[46:0] T15470;
  wire[46:0] T15471;
  wire T15472;
  wire T15473;
  wire[46:0] T15474;
  wire[46:0] T15475;
  wire[46:0] twiddle4_2_84_real;
  wire[46:0] T15476;
  wire[45:0] T15477;
  wire[45:0] T15478;
  wire T15479;
  wire[46:0] T15480;
  wire[46:0] T15481;
  wire[46:0] twiddle4_2_85_real;
  wire[46:0] T15482;
  wire[45:0] T15483;
  wire[45:0] T15484;
  wire T15485;
  wire[46:0] T15486;
  wire[46:0] T15487;
  wire T15488;
  wire[46:0] T15489;
  wire[46:0] twiddle4_2_86_real;
  wire[46:0] T15490;
  wire[46:0] T15491;
  wire[46:0] T15492;
  wire[46:0] T15493;
  wire[46:0] twiddle4_2_87_real;
  wire[46:0] T15494;
  wire[46:0] T15495;
  wire[46:0] T15496;
  wire[46:0] T15497;
  wire T15498;
  wire T15499;
  wire T15500;
  wire[46:0] T15501;
  wire[46:0] T15502;
  wire[46:0] T15503;
  wire[46:0] twiddle4_2_88_real;
  wire[46:0] T15504;
  wire[46:0] T15505;
  wire[46:0] T15506;
  wire[46:0] T15507;
  wire[46:0] twiddle4_2_89_real;
  wire[46:0] T15508;
  wire[46:0] T15509;
  wire[46:0] T15510;
  wire[46:0] T15511;
  wire T15512;
  wire[46:0] T15513;
  wire[46:0] twiddle4_2_90_real;
  wire[46:0] T15514;
  wire[46:0] T15515;
  wire[46:0] T15516;
  wire[46:0] T15517;
  wire[46:0] twiddle4_2_91_real;
  wire[46:0] T15518;
  wire[46:0] T15519;
  wire[46:0] T15520;
  wire[46:0] T15521;
  wire T15522;
  wire T15523;
  wire[46:0] T15524;
  wire[46:0] T15525;
  wire[46:0] twiddle4_2_92_real;
  wire[46:0] T15526;
  wire[46:0] T15527;
  wire[46:0] T15528;
  wire[46:0] T15529;
  wire[46:0] twiddle4_2_93_real;
  wire[46:0] T15530;
  wire[46:0] T15531;
  wire[46:0] T15532;
  wire[46:0] T15533;
  wire T15534;
  wire[46:0] T15535;
  wire[46:0] twiddle4_2_94_real;
  wire[46:0] T15536;
  wire[46:0] T15537;
  wire[46:0] T15538;
  wire[46:0] T15539;
  wire[46:0] twiddle4_2_95_real;
  wire[46:0] T15540;
  wire[46:0] T15541;
  wire[46:0] T15542;
  wire[46:0] T15543;
  wire T15544;
  wire T15545;
  wire T15546;
  wire T15547;
  wire T15548;
  wire[46:0] T15549;
  wire[46:0] T15550;
  wire[46:0] T15551;
  wire[46:0] T15552;
  wire[46:0] T15553;
  wire[46:0] twiddle4_2_96_real;
  wire[46:0] T15554;
  wire[46:0] T15555;
  wire[46:0] T15556;
  wire[46:0] T15557;
  wire[46:0] twiddle4_2_97_real;
  wire[46:0] T15558;
  wire[46:0] T15559;
  wire[46:0] T15560;
  wire[46:0] T15561;
  wire T15562;
  wire[46:0] T15563;
  wire[46:0] twiddle4_2_98_real;
  wire[46:0] T15564;
  wire[46:0] T15565;
  wire[46:0] T15566;
  wire[46:0] T15567;
  wire[46:0] twiddle4_2_99_real;
  wire[46:0] T15568;
  wire[46:0] T15569;
  wire[46:0] T15570;
  wire[46:0] T15571;
  wire T15572;
  wire T15573;
  wire[46:0] T15574;
  wire[46:0] T15575;
  wire[46:0] twiddle4_2_100_real;
  wire[46:0] T15576;
  wire[46:0] T15577;
  wire[46:0] T15578;
  wire[46:0] T15579;
  wire[46:0] twiddle4_2_101_real;
  wire[46:0] T15580;
  wire[46:0] T15581;
  wire[46:0] T15582;
  wire[46:0] T15583;
  wire T15584;
  wire[46:0] T15585;
  wire[46:0] twiddle4_2_102_real;
  wire[46:0] T15586;
  wire[46:0] T15587;
  wire[46:0] T15588;
  wire[46:0] T15589;
  wire[46:0] twiddle4_2_103_real;
  wire[46:0] T15590;
  wire[46:0] T15591;
  wire[46:0] T15592;
  wire[46:0] T15593;
  wire T15594;
  wire T15595;
  wire T15596;
  wire[46:0] T15597;
  wire[46:0] T15598;
  wire[46:0] T15599;
  wire[46:0] twiddle4_2_104_real;
  wire[46:0] T15600;
  wire[46:0] T15601;
  wire[46:0] T15602;
  wire[46:0] T15603;
  wire[46:0] twiddle4_2_105_real;
  wire[46:0] T15604;
  wire[46:0] T15605;
  wire[46:0] T15606;
  wire[46:0] T15607;
  wire T15608;
  wire[46:0] T15609;
  wire[46:0] twiddle4_2_106_real;
  wire[46:0] T15610;
  wire[46:0] T15611;
  wire[46:0] T15612;
  wire[46:0] T15613;
  wire[46:0] twiddle4_2_107_real;
  wire[46:0] T15614;
  wire[46:0] T15615;
  wire[46:0] T15616;
  wire[46:0] T15617;
  wire T15618;
  wire T15619;
  wire[46:0] T15620;
  wire[46:0] T15621;
  wire[46:0] twiddle4_2_108_real;
  wire[46:0] T15622;
  wire[46:0] T15623;
  wire[46:0] T15624;
  wire[46:0] T15625;
  wire[46:0] twiddle4_2_109_real;
  wire[46:0] T15626;
  wire[46:0] T15627;
  wire[46:0] T15628;
  wire[46:0] T15629;
  wire T15630;
  wire[46:0] T15631;
  wire[46:0] twiddle4_2_110_real;
  wire[46:0] T15632;
  wire[46:0] T15633;
  wire[46:0] T15634;
  wire[46:0] T15635;
  wire[46:0] twiddle4_2_111_real;
  wire[46:0] T15636;
  wire[46:0] T15637;
  wire[46:0] T15638;
  wire[46:0] T15639;
  wire T15640;
  wire T15641;
  wire T15642;
  wire T15643;
  wire[46:0] T15644;
  wire[46:0] T15645;
  wire[46:0] T15646;
  wire[46:0] T15647;
  wire[46:0] twiddle4_2_112_real;
  wire[46:0] T15648;
  wire[46:0] T15649;
  wire[46:0] T15650;
  wire[46:0] T15651;
  wire[46:0] twiddle4_2_113_real;
  wire[46:0] T15652;
  wire[46:0] T15653;
  wire[46:0] T15654;
  wire[46:0] T15655;
  wire T15656;
  wire[46:0] T15657;
  wire[46:0] twiddle4_2_114_real;
  wire[46:0] T15658;
  wire[46:0] T15659;
  wire[46:0] T15660;
  wire[46:0] T15661;
  wire[46:0] twiddle4_2_115_real;
  wire[46:0] T15662;
  wire[46:0] T15663;
  wire[46:0] T15664;
  wire[46:0] T15665;
  wire T15666;
  wire T15667;
  wire[46:0] T15668;
  wire[46:0] T15669;
  wire[46:0] twiddle4_2_116_real;
  wire[46:0] T15670;
  wire[46:0] T15671;
  wire[46:0] T15672;
  wire[46:0] T15673;
  wire[46:0] twiddle4_2_117_real;
  wire[46:0] T15674;
  wire[46:0] T15675;
  wire[46:0] T15676;
  wire[46:0] T15677;
  wire T15678;
  wire[46:0] T15679;
  wire[46:0] twiddle4_2_118_real;
  wire[46:0] T15680;
  wire[46:0] T15681;
  wire[46:0] T15682;
  wire[46:0] T15683;
  wire[46:0] twiddle4_2_119_real;
  wire[46:0] T15684;
  wire[46:0] T15685;
  wire[46:0] T15686;
  wire[46:0] T15687;
  wire T15688;
  wire T15689;
  wire T15690;
  wire[46:0] T15691;
  wire[46:0] T15692;
  wire[46:0] T15693;
  wire[46:0] twiddle4_2_120_real;
  wire[46:0] T15694;
  wire[46:0] T15695;
  wire[46:0] T15696;
  wire[46:0] T15697;
  wire[46:0] twiddle4_2_121_real;
  wire[46:0] T15698;
  wire[46:0] T15699;
  wire[46:0] T15700;
  wire[46:0] T15701;
  wire T15702;
  wire[46:0] T15703;
  wire[46:0] twiddle4_2_122_real;
  wire[46:0] T15704;
  wire[46:0] T15705;
  wire[46:0] T15706;
  wire[46:0] T15707;
  wire[46:0] twiddle4_2_123_real;
  wire[46:0] T15708;
  wire[46:0] T15709;
  wire[46:0] T15710;
  wire[46:0] T15711;
  wire T15712;
  wire T15713;
  wire[46:0] T15714;
  wire[46:0] T15715;
  wire[46:0] twiddle4_2_124_real;
  wire[46:0] T15716;
  wire[46:0] T15717;
  wire[46:0] T15718;
  wire[46:0] T15719;
  wire[46:0] twiddle4_2_125_real;
  wire[46:0] T15720;
  wire[46:0] T15721;
  wire[46:0] T15722;
  wire[46:0] T15723;
  wire T15724;
  wire[46:0] T15725;
  wire[46:0] twiddle4_2_126_real;
  wire[46:0] T15726;
  wire[46:0] T15727;
  wire[46:0] T15728;
  wire[46:0] T15729;
  wire[46:0] twiddle4_2_127_real;
  wire[46:0] T15730;
  wire[46:0] T15731;
  wire[46:0] T15732;
  wire[46:0] T15733;
  wire T15734;
  wire T15735;
  wire T15736;
  wire T15737;
  wire T15738;
  wire T15739;
  wire T15740;
  wire T15741;
  wire[47:0] T15742;
  wire[46:0] T15743;
  wire[46:0] T15744;
  wire[46:0] T15745;
  wire[46:0] T15746;
  wire[46:0] T15747;
  wire[46:0] T15748;
  wire[46:0] T15749;
  wire[46:0] twiddle4_2_128_real;
  wire[46:0] T15750;
  wire[46:0] T15751;
  wire[46:0] T15752;
  wire[46:0] T15753;
  wire[46:0] twiddle4_2_129_real;
  wire[46:0] T15754;
  wire[46:0] T15755;
  wire[46:0] T15756;
  wire[46:0] T15757;
  wire T15758;
  wire[46:0] T15759;
  wire[46:0] twiddle4_2_130_real;
  wire[46:0] T15760;
  wire[46:0] T15761;
  wire[46:0] T15762;
  wire[46:0] T15763;
  wire[46:0] twiddle4_2_131_real;
  wire[46:0] T15764;
  wire[46:0] T15765;
  wire[46:0] T15766;
  wire[46:0] T15767;
  wire T15768;
  wire T15769;
  wire[46:0] T15770;
  wire[46:0] T15771;
  wire[46:0] twiddle4_2_132_real;
  wire[46:0] T15772;
  wire[46:0] T15773;
  wire[46:0] T15774;
  wire[46:0] T15775;
  wire[46:0] twiddle4_2_133_real;
  wire[46:0] T15776;
  wire[46:0] T15777;
  wire[46:0] T15778;
  wire[46:0] T15779;
  wire T15780;
  wire[46:0] T15781;
  wire[46:0] twiddle4_2_134_real;
  wire[46:0] T15782;
  wire[46:0] T15783;
  wire[46:0] T15784;
  wire[46:0] T15785;
  wire[46:0] twiddle4_2_135_real;
  wire[46:0] T15786;
  wire[46:0] T15787;
  wire[46:0] T15788;
  wire[46:0] T15789;
  wire T15790;
  wire T15791;
  wire T15792;
  wire[46:0] T15793;
  wire[46:0] T15794;
  wire[46:0] T15795;
  wire[46:0] twiddle4_2_136_real;
  wire[46:0] T15796;
  wire[46:0] T15797;
  wire[46:0] T15798;
  wire[46:0] T15799;
  wire[46:0] twiddle4_2_137_real;
  wire[46:0] T15800;
  wire[46:0] T15801;
  wire[46:0] T15802;
  wire[46:0] T15803;
  wire T15804;
  wire[46:0] T15805;
  wire[46:0] twiddle4_2_138_real;
  wire[46:0] T15806;
  wire[46:0] T15807;
  wire[46:0] T15808;
  wire[46:0] T15809;
  wire[46:0] twiddle4_2_139_real;
  wire[46:0] T15810;
  wire[46:0] T15811;
  wire[46:0] T15812;
  wire[46:0] T15813;
  wire T15814;
  wire T15815;
  wire[46:0] T15816;
  wire[46:0] T15817;
  wire[46:0] twiddle4_2_140_real;
  wire[46:0] T15818;
  wire[46:0] T15819;
  wire[46:0] T15820;
  wire[46:0] T15821;
  wire[46:0] twiddle4_2_141_real;
  wire[46:0] T15822;
  wire[46:0] T15823;
  wire[46:0] T15824;
  wire[46:0] T15825;
  wire T15826;
  wire[46:0] T15827;
  wire[46:0] twiddle4_2_142_real;
  wire[46:0] T15828;
  wire[46:0] T15829;
  wire[46:0] T15830;
  wire[46:0] T15831;
  wire[46:0] twiddle4_2_143_real;
  wire[46:0] T15832;
  wire[46:0] T15833;
  wire[46:0] T15834;
  wire[46:0] T15835;
  wire T15836;
  wire T15837;
  wire T15838;
  wire T15839;
  wire[46:0] T15840;
  wire[46:0] T15841;
  wire[46:0] T15842;
  wire[46:0] T15843;
  wire[46:0] twiddle4_2_144_real;
  wire[46:0] T15844;
  wire[46:0] T15845;
  wire[46:0] T15846;
  wire[46:0] T15847;
  wire[46:0] twiddle4_2_145_real;
  wire[46:0] T15848;
  wire[46:0] T15849;
  wire[46:0] T15850;
  wire[46:0] T15851;
  wire T15852;
  wire[46:0] T15853;
  wire[46:0] twiddle4_2_146_real;
  wire[46:0] T15854;
  wire[46:0] T15855;
  wire[46:0] T15856;
  wire[46:0] T15857;
  wire[46:0] twiddle4_2_147_real;
  wire[46:0] T15858;
  wire[46:0] T15859;
  wire[46:0] T15860;
  wire[46:0] T15861;
  wire T15862;
  wire T15863;
  wire[46:0] T15864;
  wire[46:0] T15865;
  wire[46:0] twiddle4_2_148_real;
  wire[46:0] T15866;
  wire[46:0] T15867;
  wire[46:0] T15868;
  wire[46:0] T15869;
  wire[46:0] twiddle4_2_149_real;
  wire[46:0] T15870;
  wire[46:0] T15871;
  wire[46:0] T15872;
  wire[46:0] T15873;
  wire T15874;
  wire[46:0] T15875;
  wire[46:0] twiddle4_2_150_real;
  wire[46:0] T15876;
  wire[46:0] T15877;
  wire[46:0] T15878;
  wire[46:0] T15879;
  wire[46:0] twiddle4_2_151_real;
  wire[46:0] T15880;
  wire[46:0] T15881;
  wire[46:0] T15882;
  wire[46:0] T15883;
  wire T15884;
  wire T15885;
  wire T15886;
  wire[46:0] T15887;
  wire[46:0] T15888;
  wire[46:0] T15889;
  wire[46:0] twiddle4_2_152_real;
  wire[46:0] T15890;
  wire[46:0] T15891;
  wire[46:0] T15892;
  wire[46:0] T15893;
  wire[46:0] twiddle4_2_153_real;
  wire[46:0] T15894;
  wire[46:0] T15895;
  wire[46:0] T15896;
  wire[46:0] T15897;
  wire T15898;
  wire[46:0] T15899;
  wire[46:0] twiddle4_2_154_real;
  wire[46:0] T15900;
  wire[46:0] T15901;
  wire[46:0] T15902;
  wire[46:0] T15903;
  wire[46:0] twiddle4_2_155_real;
  wire[46:0] T15904;
  wire[46:0] T15905;
  wire[46:0] T15906;
  wire[46:0] T15907;
  wire T15908;
  wire T15909;
  wire[46:0] T15910;
  wire[46:0] T15911;
  wire[46:0] twiddle4_2_156_real;
  wire[46:0] T15912;
  wire[46:0] T15913;
  wire[46:0] T15914;
  wire[46:0] T15915;
  wire[46:0] twiddle4_2_157_real;
  wire[46:0] T15916;
  wire[46:0] T15917;
  wire[46:0] T15918;
  wire[46:0] T15919;
  wire T15920;
  wire[46:0] T15921;
  wire[46:0] twiddle4_2_158_real;
  wire[46:0] T15922;
  wire[46:0] T15923;
  wire[46:0] T15924;
  wire[46:0] T15925;
  wire[46:0] twiddle4_2_159_real;
  wire[46:0] T15926;
  wire[46:0] T15927;
  wire[46:0] T15928;
  wire[46:0] T15929;
  wire T15930;
  wire T15931;
  wire T15932;
  wire T15933;
  wire T15934;
  wire[46:0] T15935;
  wire[46:0] T15936;
  wire[46:0] T15937;
  wire[46:0] T15938;
  wire[46:0] T15939;
  wire[46:0] twiddle4_2_160_real;
  wire[46:0] T15940;
  wire[46:0] T15941;
  wire[46:0] T15942;
  wire[46:0] T15943;
  wire[46:0] twiddle4_2_161_real;
  wire[46:0] T15944;
  wire[46:0] T15945;
  wire[46:0] T15946;
  wire[46:0] T15947;
  wire T15948;
  wire[46:0] T15949;
  wire[46:0] twiddle4_2_162_real;
  wire[46:0] T15950;
  wire[46:0] T15951;
  wire[46:0] T15952;
  wire[46:0] T15953;
  wire[46:0] twiddle4_2_163_real;
  wire[46:0] T15954;
  wire[46:0] T15955;
  wire[46:0] T15956;
  wire[46:0] T15957;
  wire T15958;
  wire T15959;
  wire[46:0] T15960;
  wire[46:0] T15961;
  wire[46:0] twiddle4_2_164_real;
  wire[46:0] T15962;
  wire[46:0] T15963;
  wire[46:0] T15964;
  wire[46:0] T15965;
  wire[46:0] twiddle4_2_165_real;
  wire[46:0] T15966;
  wire[46:0] T15967;
  wire[46:0] T15968;
  wire[46:0] T15969;
  wire T15970;
  wire[46:0] T15971;
  wire[46:0] twiddle4_2_166_real;
  wire[46:0] T15972;
  wire[46:0] T15973;
  wire[46:0] T15974;
  wire[46:0] T15975;
  wire[46:0] twiddle4_2_167_real;
  wire[46:0] T15976;
  wire[46:0] T15977;
  wire[46:0] T15978;
  wire[46:0] T15979;
  wire T15980;
  wire T15981;
  wire T15982;
  wire[46:0] T15983;
  wire[46:0] T15984;
  wire[46:0] T15985;
  wire[46:0] twiddle4_2_168_real;
  wire[46:0] T15986;
  wire[46:0] T15987;
  wire[46:0] T15988;
  wire[46:0] T15989;
  wire[46:0] twiddle4_2_169_real;
  wire[46:0] T15990;
  wire[46:0] T15991;
  wire[46:0] T15992;
  wire[46:0] T15993;
  wire T15994;
  wire[46:0] T15995;
  wire[46:0] twiddle4_2_170_real;
  wire[46:0] T15996;
  wire[46:0] T15997;
  wire[46:0] T15998;
  wire[46:0] T15999;
  wire[46:0] twiddle4_2_171_real;
  wire[46:0] T16000;
  wire[46:0] T16001;
  wire[46:0] T16002;
  wire[45:0] T16003;
  wire[45:0] T16004;
  wire T16005;
  wire T16006;
  wire T16007;
  wire[46:0] T16008;
  wire[46:0] T16009;
  wire[46:0] twiddle4_2_172_real;
  wire[46:0] T16010;
  wire[46:0] T16011;
  wire[46:0] T16012;
  wire[45:0] T16013;
  wire[45:0] T16014;
  wire T16015;
  wire[46:0] twiddle4_2_173_real;
  wire[46:0] T16016;
  wire[46:0] T16017;
  wire[46:0] T16018;
  wire[45:0] T16019;
  wire[45:0] T16020;
  wire T16021;
  wire T16022;
  wire[46:0] T16023;
  wire[46:0] twiddle4_2_174_real;
  wire[46:0] T16024;
  wire[46:0] T16025;
  wire[46:0] T16026;
  wire[45:0] T16027;
  wire[45:0] T16028;
  wire T16029;
  wire[46:0] twiddle4_2_175_real;
  wire[46:0] T16030;
  wire[46:0] T16031;
  wire[46:0] T16032;
  wire[45:0] T16033;
  wire[45:0] T16034;
  wire T16035;
  wire T16036;
  wire T16037;
  wire T16038;
  wire T16039;
  wire[46:0] T16040;
  wire[46:0] T16041;
  wire[46:0] T16042;
  wire[46:0] T16043;
  wire[46:0] twiddle4_2_176_real;
  wire[46:0] T16044;
  wire[46:0] T16045;
  wire[46:0] T16046;
  wire[45:0] T16047;
  wire[45:0] T16048;
  wire T16049;
  wire[46:0] twiddle4_2_177_real;
  wire[46:0] T16050;
  wire[46:0] T16051;
  wire[46:0] T16052;
  wire[45:0] T16053;
  wire[45:0] T16054;
  wire T16055;
  wire T16056;
  wire[46:0] T16057;
  wire[46:0] twiddle4_2_178_real;
  wire[46:0] T16058;
  wire[46:0] T16059;
  wire[46:0] T16060;
  wire[45:0] T16061;
  wire[45:0] T16062;
  wire T16063;
  wire[46:0] twiddle4_2_179_real;
  wire[46:0] T16064;
  wire[46:0] T16065;
  wire[46:0] T16066;
  wire[45:0] T16067;
  wire[45:0] T16068;
  wire T16069;
  wire T16070;
  wire T16071;
  wire[46:0] T16072;
  wire[46:0] T16073;
  wire[46:0] twiddle4_2_180_real;
  wire[46:0] T16074;
  wire[46:0] T16075;
  wire[46:0] T16076;
  wire[45:0] T16077;
  wire[45:0] T16078;
  wire T16079;
  wire[46:0] twiddle4_2_181_real;
  wire[46:0] T16080;
  wire[46:0] T16081;
  wire[46:0] T16082;
  wire[45:0] T16083;
  wire[45:0] T16084;
  wire T16085;
  wire T16086;
  wire[46:0] T16087;
  wire[46:0] twiddle4_2_182_real;
  wire[46:0] T16088;
  wire[46:0] T16089;
  wire[46:0] T16090;
  wire[45:0] T16091;
  wire[45:0] T16092;
  wire T16093;
  wire[46:0] twiddle4_2_183_real;
  wire[46:0] T16094;
  wire[46:0] T16095;
  wire[46:0] T16096;
  wire[45:0] T16097;
  wire[45:0] T16098;
  wire T16099;
  wire T16100;
  wire T16101;
  wire T16102;
  wire[46:0] T16103;
  wire[46:0] T16104;
  wire[46:0] T16105;
  wire[46:0] twiddle4_2_184_real;
  wire[46:0] T16106;
  wire[46:0] T16107;
  wire[46:0] T16108;
  wire[45:0] T16109;
  wire[45:0] T16110;
  wire T16111;
  wire[46:0] twiddle4_2_185_real;
  wire[46:0] T16112;
  wire[46:0] T16113;
  wire[46:0] T16114;
  wire[45:0] T16115;
  wire[45:0] T16116;
  wire T16117;
  wire T16118;
  wire[46:0] T16119;
  wire[46:0] twiddle4_2_186_real;
  wire[46:0] T16120;
  wire[46:0] T16121;
  wire[46:0] T16122;
  wire[45:0] T16123;
  wire[45:0] T16124;
  wire T16125;
  wire[46:0] twiddle4_2_187_real;
  wire[46:0] T16126;
  wire[46:0] T16127;
  wire[46:0] T16128;
  wire[45:0] T16129;
  wire[45:0] T16130;
  wire T16131;
  wire T16132;
  wire T16133;
  wire[46:0] T16134;
  wire[46:0] T16135;
  wire[46:0] twiddle4_2_188_real;
  wire[46:0] T16136;
  wire[46:0] T16137;
  wire[46:0] T16138;
  wire[45:0] T16139;
  wire[45:0] T16140;
  wire T16141;
  wire[46:0] twiddle4_2_189_real;
  wire[46:0] T16142;
  wire[46:0] T16143;
  wire[46:0] T16144;
  wire[45:0] T16145;
  wire[45:0] T16146;
  wire T16147;
  wire T16148;
  wire[46:0] T16149;
  wire[46:0] twiddle4_2_190_real;
  wire[46:0] T16150;
  wire[46:0] T16151;
  wire[46:0] T16152;
  wire[45:0] T16153;
  wire[45:0] T16154;
  wire T16155;
  wire[46:0] twiddle4_2_191_real;
  wire[46:0] T16156;
  wire[46:0] T16157;
  wire[46:0] T16158;
  wire[45:0] T16159;
  wire[45:0] T16160;
  wire T16161;
  wire T16162;
  wire T16163;
  wire T16164;
  wire T16165;
  wire T16166;
  wire T16167;
  wire[46:0] T16168;
  wire[46:0] T16169;
  wire[46:0] T16170;
  wire[46:0] T16171;
  wire[46:0] T16172;
  wire[46:0] T16173;
  wire[46:0] twiddle4_2_192_real;
  wire[46:0] T16174;
  wire[46:0] T16175;
  wire[46:0] T16176;
  wire[45:0] T16177;
  wire[45:0] T16178;
  wire T16179;
  wire[46:0] twiddle4_2_193_real;
  wire[46:0] T16180;
  wire[46:0] T16181;
  wire[46:0] T16182;
  wire[45:0] T16183;
  wire[45:0] T16184;
  wire T16185;
  wire T16186;
  wire[46:0] T16187;
  wire[46:0] twiddle4_2_194_real;
  wire[46:0] T16188;
  wire[46:0] T16189;
  wire[46:0] T16190;
  wire[45:0] T16191;
  wire[45:0] T16192;
  wire T16193;
  wire[46:0] twiddle4_2_195_real;
  wire[46:0] T16194;
  wire[46:0] T16195;
  wire[46:0] T16196;
  wire[45:0] T16197;
  wire[45:0] T16198;
  wire T16199;
  wire T16200;
  wire T16201;
  wire[46:0] T16202;
  wire[46:0] T16203;
  wire[46:0] twiddle4_2_196_real;
  wire[46:0] T16204;
  wire[46:0] T16205;
  wire[46:0] T16206;
  wire[45:0] T16207;
  wire[45:0] T16208;
  wire T16209;
  wire[46:0] twiddle4_2_197_real;
  wire[46:0] T16210;
  wire[46:0] T16211;
  wire[46:0] T16212;
  wire[45:0] T16213;
  wire[45:0] T16214;
  wire T16215;
  wire T16216;
  wire[46:0] T16217;
  wire[46:0] twiddle4_2_198_real;
  wire[46:0] T16218;
  wire[46:0] T16219;
  wire[46:0] T16220;
  wire[45:0] T16221;
  wire[45:0] T16222;
  wire T16223;
  wire[46:0] twiddle4_2_199_real;
  wire[46:0] T16224;
  wire[46:0] T16225;
  wire[46:0] T16226;
  wire[45:0] T16227;
  wire[45:0] T16228;
  wire T16229;
  wire T16230;
  wire T16231;
  wire T16232;
  wire[46:0] T16233;
  wire[46:0] T16234;
  wire[46:0] T16235;
  wire[46:0] twiddle4_2_200_real;
  wire[46:0] T16236;
  wire[46:0] T16237;
  wire[46:0] T16238;
  wire[45:0] T16239;
  wire[45:0] T16240;
  wire T16241;
  wire[46:0] twiddle4_2_201_real;
  wire[46:0] T16242;
  wire[46:0] T16243;
  wire[46:0] T16244;
  wire[45:0] T16245;
  wire[45:0] T16246;
  wire T16247;
  wire T16248;
  wire[46:0] T16249;
  wire[46:0] twiddle4_2_202_real;
  wire[46:0] T16250;
  wire[46:0] T16251;
  wire[46:0] T16252;
  wire[45:0] T16253;
  wire[45:0] T16254;
  wire T16255;
  wire[46:0] twiddle4_2_203_real;
  wire[46:0] T16256;
  wire[46:0] T16257;
  wire[46:0] T16258;
  wire[45:0] T16259;
  wire[45:0] T16260;
  wire T16261;
  wire T16262;
  wire T16263;
  wire[46:0] T16264;
  wire[46:0] T16265;
  wire[46:0] twiddle4_2_204_real;
  wire[46:0] T16266;
  wire[46:0] T16267;
  wire[46:0] T16268;
  wire[45:0] T16269;
  wire[45:0] T16270;
  wire T16271;
  wire[46:0] twiddle4_2_205_real;
  wire[46:0] T16272;
  wire[46:0] T16273;
  wire[46:0] T16274;
  wire[45:0] T16275;
  wire[45:0] T16276;
  wire T16277;
  wire T16278;
  wire[46:0] T16279;
  wire[46:0] twiddle4_2_206_real;
  wire[46:0] T16280;
  wire[46:0] T16281;
  wire[46:0] T16282;
  wire[45:0] T16283;
  wire[45:0] T16284;
  wire T16285;
  wire[46:0] twiddle4_2_207_real;
  wire[46:0] T16286;
  wire[46:0] T16287;
  wire[46:0] T16288;
  wire[45:0] T16289;
  wire[45:0] T16290;
  wire T16291;
  wire T16292;
  wire T16293;
  wire T16294;
  wire T16295;
  wire[46:0] T16296;
  wire[46:0] T16297;
  wire[46:0] T16298;
  wire[46:0] T16299;
  wire[46:0] twiddle4_2_208_real;
  wire[46:0] T16300;
  wire[46:0] T16301;
  wire[46:0] T16302;
  wire[45:0] T16303;
  wire[45:0] T16304;
  wire T16305;
  wire[46:0] twiddle4_2_209_real;
  wire[46:0] T16306;
  wire[46:0] T16307;
  wire[46:0] T16308;
  wire[45:0] T16309;
  wire[45:0] T16310;
  wire T16311;
  wire T16312;
  wire[46:0] T16313;
  wire[46:0] twiddle4_2_210_real;
  wire[46:0] T16314;
  wire[46:0] T16315;
  wire[46:0] T16316;
  wire[45:0] T16317;
  wire[45:0] T16318;
  wire T16319;
  wire[46:0] twiddle4_2_211_real;
  wire[46:0] T16320;
  wire[46:0] T16321;
  wire[46:0] T16322;
  wire[45:0] T16323;
  wire[45:0] T16324;
  wire T16325;
  wire T16326;
  wire T16327;
  wire[46:0] T16328;
  wire[46:0] T16329;
  wire[46:0] twiddle4_2_212_real;
  wire[46:0] T16330;
  wire[46:0] T16331;
  wire[46:0] T16332;
  wire[45:0] T16333;
  wire[45:0] T16334;
  wire T16335;
  wire[46:0] twiddle4_2_213_real;
  wire[46:0] T16336;
  wire[46:0] T16337;
  wire[46:0] T16338;
  wire[45:0] T16339;
  wire[45:0] T16340;
  wire T16341;
  wire T16342;
  wire[46:0] T16343;
  wire[46:0] twiddle4_2_214_real;
  wire[46:0] T16344;
  wire[46:0] T16345;
  wire[46:0] T16346;
  wire[45:0] T16347;
  wire[45:0] T16348;
  wire T16349;
  wire[46:0] twiddle4_2_215_real;
  wire[46:0] T16350;
  wire[46:0] T16351;
  wire[46:0] T16352;
  wire[44:0] T16353;
  wire[44:0] T16354;
  wire[1:0] T16355;
  wire T16356;
  wire T16357;
  wire T16358;
  wire T16359;
  wire[46:0] T16360;
  wire[46:0] T16361;
  wire[46:0] T16362;
  wire[46:0] twiddle4_2_216_real;
  wire[46:0] T16363;
  wire[46:0] T16364;
  wire[46:0] T16365;
  wire[44:0] T16366;
  wire[44:0] T16367;
  wire[1:0] T16368;
  wire T16369;
  wire[46:0] twiddle4_2_217_real;
  wire[46:0] T16370;
  wire[46:0] T16371;
  wire[46:0] T16372;
  wire[44:0] T16373;
  wire[44:0] T16374;
  wire[1:0] T16375;
  wire T16376;
  wire T16377;
  wire[46:0] T16378;
  wire[46:0] twiddle4_2_218_real;
  wire[46:0] T16379;
  wire[46:0] T16380;
  wire[46:0] T16381;
  wire[44:0] T16382;
  wire[44:0] T16383;
  wire[1:0] T16384;
  wire T16385;
  wire[46:0] twiddle4_2_219_real;
  wire[46:0] T16386;
  wire[46:0] T16387;
  wire[46:0] T16388;
  wire[44:0] T16389;
  wire[44:0] T16390;
  wire[1:0] T16391;
  wire T16392;
  wire T16393;
  wire T16394;
  wire[46:0] T16395;
  wire[46:0] T16396;
  wire[46:0] twiddle4_2_220_real;
  wire[46:0] T16397;
  wire[46:0] T16398;
  wire[46:0] T16399;
  wire[44:0] T16400;
  wire[44:0] T16401;
  wire[1:0] T16402;
  wire T16403;
  wire[46:0] twiddle4_2_221_real;
  wire[46:0] T16404;
  wire[46:0] T16405;
  wire[46:0] T16406;
  wire[44:0] T16407;
  wire[44:0] T16408;
  wire[1:0] T16409;
  wire T16410;
  wire T16411;
  wire[46:0] T16412;
  wire[46:0] twiddle4_2_222_real;
  wire[46:0] T16413;
  wire[46:0] T16414;
  wire[46:0] T16415;
  wire[44:0] T16416;
  wire[44:0] T16417;
  wire[1:0] T16418;
  wire T16419;
  wire[46:0] twiddle4_2_223_real;
  wire[46:0] T16420;
  wire[46:0] T16421;
  wire[46:0] T16422;
  wire[44:0] T16423;
  wire[44:0] T16424;
  wire[1:0] T16425;
  wire T16426;
  wire T16427;
  wire T16428;
  wire T16429;
  wire T16430;
  wire T16431;
  wire[46:0] T16432;
  wire[46:0] T16433;
  wire[46:0] T16434;
  wire[46:0] T16435;
  wire[46:0] T16436;
  wire[46:0] twiddle4_2_224_real;
  wire[46:0] T16437;
  wire[46:0] T16438;
  wire[46:0] T16439;
  wire[44:0] T16440;
  wire[44:0] T16441;
  wire[1:0] T16442;
  wire T16443;
  wire[46:0] twiddle4_2_225_real;
  wire[46:0] T16444;
  wire[46:0] T16445;
  wire[46:0] T16446;
  wire[44:0] T16447;
  wire[44:0] T16448;
  wire[1:0] T16449;
  wire T16450;
  wire T16451;
  wire[46:0] T16452;
  wire[46:0] twiddle4_2_226_real;
  wire[46:0] T16453;
  wire[46:0] T16454;
  wire[46:0] T16455;
  wire[44:0] T16456;
  wire[44:0] T16457;
  wire[1:0] T16458;
  wire T16459;
  wire[46:0] twiddle4_2_227_real;
  wire[46:0] T16460;
  wire[46:0] T16461;
  wire[46:0] T16462;
  wire[44:0] T16463;
  wire[44:0] T16464;
  wire[1:0] T16465;
  wire T16466;
  wire T16467;
  wire T16468;
  wire[46:0] T16469;
  wire[46:0] T16470;
  wire[46:0] twiddle4_2_228_real;
  wire[46:0] T16471;
  wire[46:0] T16472;
  wire[46:0] T16473;
  wire[44:0] T16474;
  wire[44:0] T16475;
  wire[1:0] T16476;
  wire T16477;
  wire[46:0] twiddle4_2_229_real;
  wire[46:0] T16478;
  wire[46:0] T16479;
  wire[46:0] T16480;
  wire[44:0] T16481;
  wire[44:0] T16482;
  wire[1:0] T16483;
  wire T16484;
  wire T16485;
  wire[46:0] T16486;
  wire[46:0] twiddle4_2_230_real;
  wire[46:0] T16487;
  wire[46:0] T16488;
  wire[46:0] T16489;
  wire[44:0] T16490;
  wire[44:0] T16491;
  wire[1:0] T16492;
  wire T16493;
  wire[46:0] twiddle4_2_231_real;
  wire[46:0] T16494;
  wire[46:0] T16495;
  wire[46:0] T16496;
  wire[44:0] T16497;
  wire[44:0] T16498;
  wire[1:0] T16499;
  wire T16500;
  wire T16501;
  wire T16502;
  wire T16503;
  wire[46:0] T16504;
  wire[46:0] T16505;
  wire[46:0] T16506;
  wire[46:0] twiddle4_2_232_real;
  wire[46:0] T16507;
  wire[46:0] T16508;
  wire[46:0] T16509;
  wire[44:0] T16510;
  wire[44:0] T16511;
  wire[1:0] T16512;
  wire T16513;
  wire[46:0] twiddle4_2_233_real;
  wire[46:0] T16514;
  wire[46:0] T16515;
  wire[46:0] T16516;
  wire[44:0] T16517;
  wire[44:0] T16518;
  wire[1:0] T16519;
  wire T16520;
  wire T16521;
  wire[46:0] T16522;
  wire[46:0] twiddle4_2_234_real;
  wire[46:0] T16523;
  wire[46:0] T16524;
  wire[46:0] T16525;
  wire[44:0] T16526;
  wire[44:0] T16527;
  wire[1:0] T16528;
  wire T16529;
  wire[46:0] twiddle4_2_235_real;
  wire[46:0] T16530;
  wire[46:0] T16531;
  wire[46:0] T16532;
  wire[44:0] T16533;
  wire[44:0] T16534;
  wire[1:0] T16535;
  wire T16536;
  wire T16537;
  wire T16538;
  wire[46:0] T16539;
  wire[46:0] T16540;
  wire[46:0] twiddle4_2_236_real;
  wire[46:0] T16541;
  wire[46:0] T16542;
  wire[46:0] T16543;
  wire[43:0] T16544;
  wire[43:0] T16545;
  wire[2:0] T16546;
  wire T16547;
  wire[46:0] twiddle4_2_237_real;
  wire[46:0] T16548;
  wire[46:0] T16549;
  wire[46:0] T16550;
  wire[43:0] T16551;
  wire[43:0] T16552;
  wire[2:0] T16553;
  wire T16554;
  wire T16555;
  wire[46:0] T16556;
  wire[46:0] twiddle4_2_238_real;
  wire[46:0] T16557;
  wire[46:0] T16558;
  wire[46:0] T16559;
  wire[43:0] T16560;
  wire[43:0] T16561;
  wire[2:0] T16562;
  wire T16563;
  wire[46:0] twiddle4_2_239_real;
  wire[46:0] T16564;
  wire[46:0] T16565;
  wire[46:0] T16566;
  wire[43:0] T16567;
  wire[43:0] T16568;
  wire[2:0] T16569;
  wire T16570;
  wire T16571;
  wire T16572;
  wire T16573;
  wire T16574;
  wire[46:0] T16575;
  wire[46:0] T16576;
  wire[46:0] T16577;
  wire[46:0] T16578;
  wire[46:0] twiddle4_2_240_real;
  wire[46:0] T16579;
  wire[46:0] T16580;
  wire[46:0] T16581;
  wire[43:0] T16582;
  wire[43:0] T16583;
  wire[2:0] T16584;
  wire T16585;
  wire[46:0] twiddle4_2_241_real;
  wire[46:0] T16586;
  wire[46:0] T16587;
  wire[46:0] T16588;
  wire[43:0] T16589;
  wire[43:0] T16590;
  wire[2:0] T16591;
  wire T16592;
  wire T16593;
  wire[46:0] T16594;
  wire[46:0] twiddle4_2_242_real;
  wire[46:0] T16595;
  wire[46:0] T16596;
  wire[46:0] T16597;
  wire[43:0] T16598;
  wire[43:0] T16599;
  wire[2:0] T16600;
  wire T16601;
  wire[46:0] twiddle4_2_243_real;
  wire[46:0] T16602;
  wire[46:0] T16603;
  wire[46:0] T16604;
  wire[43:0] T16605;
  wire[43:0] T16606;
  wire[2:0] T16607;
  wire T16608;
  wire T16609;
  wire T16610;
  wire[46:0] T16611;
  wire[46:0] T16612;
  wire[46:0] twiddle4_2_244_real;
  wire[46:0] T16613;
  wire[46:0] T16614;
  wire[46:0] T16615;
  wire[43:0] T16616;
  wire[43:0] T16617;
  wire[2:0] T16618;
  wire T16619;
  wire[46:0] twiddle4_2_245_real;
  wire[46:0] T16620;
  wire[46:0] T16621;
  wire[46:0] T16622;
  wire[43:0] T16623;
  wire[43:0] T16624;
  wire[2:0] T16625;
  wire T16626;
  wire T16627;
  wire[46:0] T16628;
  wire[46:0] twiddle4_2_246_real;
  wire[46:0] T16629;
  wire[46:0] T16630;
  wire[46:0] T16631;
  wire[42:0] T16632;
  wire[42:0] T16633;
  wire[3:0] T16634;
  wire T16635;
  wire[46:0] twiddle4_2_247_real;
  wire[46:0] T16636;
  wire[46:0] T16637;
  wire[46:0] T16638;
  wire[42:0] T16639;
  wire[42:0] T16640;
  wire[3:0] T16641;
  wire T16642;
  wire T16643;
  wire T16644;
  wire T16645;
  wire[46:0] T16646;
  wire[46:0] T16647;
  wire[46:0] T16648;
  wire[46:0] twiddle4_2_248_real;
  wire[46:0] T16649;
  wire[46:0] T16650;
  wire[46:0] T16651;
  wire[42:0] T16652;
  wire[42:0] T16653;
  wire[3:0] T16654;
  wire T16655;
  wire[46:0] twiddle4_2_249_real;
  wire[46:0] T16656;
  wire[46:0] T16657;
  wire[46:0] T16658;
  wire[42:0] T16659;
  wire[42:0] T16660;
  wire[3:0] T16661;
  wire T16662;
  wire T16663;
  wire[46:0] T16664;
  wire[46:0] twiddle4_2_250_real;
  wire[46:0] T16665;
  wire[46:0] T16666;
  wire[46:0] T16667;
  wire[42:0] T16668;
  wire[42:0] T16669;
  wire[3:0] T16670;
  wire T16671;
  wire[46:0] twiddle4_2_251_real;
  wire[46:0] T16672;
  wire[46:0] T16673;
  wire[46:0] T16674;
  wire[41:0] T16675;
  wire[41:0] T16676;
  wire[4:0] T16677;
  wire T16678;
  wire T16679;
  wire T16680;
  wire[46:0] T16681;
  wire[46:0] T16682;
  wire[46:0] twiddle4_2_252_real;
  wire[46:0] T16683;
  wire[46:0] T16684;
  wire[46:0] T16685;
  wire[41:0] T16686;
  wire[41:0] T16687;
  wire[4:0] T16688;
  wire T16689;
  wire[46:0] twiddle4_2_253_real;
  wire[46:0] T16690;
  wire[46:0] T16691;
  wire[46:0] T16692;
  wire[41:0] T16693;
  wire[41:0] T16694;
  wire[4:0] T16695;
  wire T16696;
  wire T16697;
  wire[46:0] T16698;
  wire[46:0] twiddle4_2_254_real;
  wire[46:0] T16699;
  wire[46:0] T16700;
  wire[46:0] T16701;
  wire[40:0] T16702;
  wire[40:0] T16703;
  wire[5:0] T16704;
  wire T16705;
  wire[46:0] twiddle4_2_255_real;
  wire[46:0] T16706;
  wire[46:0] T16707;
  wire[46:0] T16708;
  wire[39:0] T16709;
  wire[39:0] T16710;
  wire[6:0] T16711;
  wire T16712;
  wire T16713;
  wire T16714;
  wire T16715;
  wire T16716;
  wire T16717;
  wire T16718;
  wire T16719;
  wire T16720;
  wire T16721;
  wire[47:0] T16722;
  wire[47:0] T16723;
  wire[47:0] T16724;
  wire[47:0] T16725;
  wire[47:0] T16726;
  wire[47:0] T16727;
  wire[47:0] T16728;
  wire[47:0] T16729;
  wire[47:0] twiddle4_2_256_real;
  wire[47:0] T16730;
  wire[47:0] T16731;
  wire[47:0] T16732;
  wire[16:0] T16733;
  wire[16:0] T16734;
  wire[30:0] T16735;
  wire T16736;
  wire[47:0] T16737;
  wire[46:0] twiddle4_2_257_real;
  wire[46:0] T16738;
  wire[46:0] T16739;
  wire[46:0] T16740;
  wire[39:0] T16741;
  wire[39:0] T16742;
  wire[6:0] T16743;
  wire T16744;
  wire T16745;
  wire T16746;
  wire[47:0] T16747;
  wire[46:0] T16748;
  wire[46:0] twiddle4_2_258_real;
  wire[46:0] T16749;
  wire[46:0] T16750;
  wire[46:0] T16751;
  wire[40:0] T16752;
  wire[40:0] T16753;
  wire[5:0] T16754;
  wire T16755;
  wire[46:0] twiddle4_2_259_real;
  wire[46:0] T16756;
  wire[46:0] T16757;
  wire[46:0] T16758;
  wire[41:0] T16759;
  wire[41:0] T16760;
  wire[4:0] T16761;
  wire T16762;
  wire T16763;
  wire T16764;
  wire T16765;
  wire[47:0] T16766;
  wire[46:0] T16767;
  wire[46:0] T16768;
  wire[46:0] twiddle4_2_260_real;
  wire[46:0] T16769;
  wire[46:0] T16770;
  wire[46:0] T16771;
  wire[41:0] T16772;
  wire[41:0] T16773;
  wire[4:0] T16774;
  wire T16775;
  wire[46:0] twiddle4_2_261_real;
  wire[46:0] T16776;
  wire[46:0] T16777;
  wire[46:0] T16778;
  wire[41:0] T16779;
  wire[41:0] T16780;
  wire[4:0] T16781;
  wire T16782;
  wire T16783;
  wire[46:0] T16784;
  wire[46:0] twiddle4_2_262_real;
  wire[46:0] T16785;
  wire[46:0] T16786;
  wire[46:0] T16787;
  wire[42:0] T16788;
  wire[42:0] T16789;
  wire[3:0] T16790;
  wire T16791;
  wire[46:0] twiddle4_2_263_real;
  wire[46:0] T16792;
  wire[46:0] T16793;
  wire[46:0] T16794;
  wire[42:0] T16795;
  wire[42:0] T16796;
  wire[3:0] T16797;
  wire T16798;
  wire T16799;
  wire T16800;
  wire T16801;
  wire T16802;
  wire[47:0] T16803;
  wire[46:0] T16804;
  wire[46:0] T16805;
  wire[46:0] T16806;
  wire[46:0] twiddle4_2_264_real;
  wire[46:0] T16807;
  wire[46:0] T16808;
  wire[46:0] T16809;
  wire[42:0] T16810;
  wire[42:0] T16811;
  wire[3:0] T16812;
  wire T16813;
  wire[46:0] twiddle4_2_265_real;
  wire[46:0] T16814;
  wire[46:0] T16815;
  wire[46:0] T16816;
  wire[42:0] T16817;
  wire[42:0] T16818;
  wire[3:0] T16819;
  wire T16820;
  wire T16821;
  wire[46:0] T16822;
  wire[46:0] twiddle4_2_266_real;
  wire[46:0] T16823;
  wire[46:0] T16824;
  wire[46:0] T16825;
  wire[42:0] T16826;
  wire[42:0] T16827;
  wire[3:0] T16828;
  wire T16829;
  wire[46:0] twiddle4_2_267_real;
  wire[46:0] T16830;
  wire[46:0] T16831;
  wire[46:0] T16832;
  wire[43:0] T16833;
  wire[43:0] T16834;
  wire[2:0] T16835;
  wire T16836;
  wire T16837;
  wire T16838;
  wire[46:0] T16839;
  wire[46:0] T16840;
  wire[46:0] twiddle4_2_268_real;
  wire[46:0] T16841;
  wire[46:0] T16842;
  wire[46:0] T16843;
  wire[43:0] T16844;
  wire[43:0] T16845;
  wire[2:0] T16846;
  wire T16847;
  wire[46:0] twiddle4_2_269_real;
  wire[46:0] T16848;
  wire[46:0] T16849;
  wire[46:0] T16850;
  wire[43:0] T16851;
  wire[43:0] T16852;
  wire[2:0] T16853;
  wire T16854;
  wire T16855;
  wire[46:0] T16856;
  wire[46:0] twiddle4_2_270_real;
  wire[46:0] T16857;
  wire[46:0] T16858;
  wire[46:0] T16859;
  wire[43:0] T16860;
  wire[43:0] T16861;
  wire[2:0] T16862;
  wire T16863;
  wire[46:0] twiddle4_2_271_real;
  wire[46:0] T16864;
  wire[46:0] T16865;
  wire[46:0] T16866;
  wire[43:0] T16867;
  wire[43:0] T16868;
  wire[2:0] T16869;
  wire T16870;
  wire T16871;
  wire T16872;
  wire T16873;
  wire T16874;
  wire T16875;
  wire[47:0] T16876;
  wire[46:0] T16877;
  wire[46:0] T16878;
  wire[46:0] T16879;
  wire[46:0] T16880;
  wire[46:0] twiddle4_2_272_real;
  wire[46:0] T16881;
  wire[46:0] T16882;
  wire[46:0] T16883;
  wire[43:0] T16884;
  wire[43:0] T16885;
  wire[2:0] T16886;
  wire T16887;
  wire[46:0] twiddle4_2_273_real;
  wire[46:0] T16888;
  wire[46:0] T16889;
  wire[46:0] T16890;
  wire[43:0] T16891;
  wire[43:0] T16892;
  wire[2:0] T16893;
  wire T16894;
  wire T16895;
  wire[46:0] T16896;
  wire[46:0] twiddle4_2_274_real;
  wire[46:0] T16897;
  wire[46:0] T16898;
  wire[46:0] T16899;
  wire[43:0] T16900;
  wire[43:0] T16901;
  wire[2:0] T16902;
  wire T16903;
  wire[46:0] twiddle4_2_275_real;
  wire[46:0] T16904;
  wire[46:0] T16905;
  wire[46:0] T16906;
  wire[43:0] T16907;
  wire[43:0] T16908;
  wire[2:0] T16909;
  wire T16910;
  wire T16911;
  wire T16912;
  wire[46:0] T16913;
  wire[46:0] T16914;
  wire[46:0] twiddle4_2_276_real;
  wire[46:0] T16915;
  wire[46:0] T16916;
  wire[46:0] T16917;
  wire[43:0] T16918;
  wire[43:0] T16919;
  wire[2:0] T16920;
  wire T16921;
  wire[46:0] twiddle4_2_277_real;
  wire[46:0] T16922;
  wire[46:0] T16923;
  wire[46:0] T16924;
  wire[44:0] T16925;
  wire[44:0] T16926;
  wire[1:0] T16927;
  wire T16928;
  wire T16929;
  wire[46:0] T16930;
  wire[46:0] twiddle4_2_278_real;
  wire[46:0] T16931;
  wire[46:0] T16932;
  wire[46:0] T16933;
  wire[44:0] T16934;
  wire[44:0] T16935;
  wire[1:0] T16936;
  wire T16937;
  wire[46:0] twiddle4_2_279_real;
  wire[46:0] T16938;
  wire[46:0] T16939;
  wire[46:0] T16940;
  wire[44:0] T16941;
  wire[44:0] T16942;
  wire[1:0] T16943;
  wire T16944;
  wire T16945;
  wire T16946;
  wire T16947;
  wire[46:0] T16948;
  wire[46:0] T16949;
  wire[46:0] T16950;
  wire[46:0] twiddle4_2_280_real;
  wire[46:0] T16951;
  wire[46:0] T16952;
  wire[46:0] T16953;
  wire[44:0] T16954;
  wire[44:0] T16955;
  wire[1:0] T16956;
  wire T16957;
  wire[46:0] twiddle4_2_281_real;
  wire[46:0] T16958;
  wire[46:0] T16959;
  wire[46:0] T16960;
  wire[44:0] T16961;
  wire[44:0] T16962;
  wire[1:0] T16963;
  wire T16964;
  wire T16965;
  wire[46:0] T16966;
  wire[46:0] twiddle4_2_282_real;
  wire[46:0] T16967;
  wire[46:0] T16968;
  wire[46:0] T16969;
  wire[44:0] T16970;
  wire[44:0] T16971;
  wire[1:0] T16972;
  wire T16973;
  wire[46:0] twiddle4_2_283_real;
  wire[46:0] T16974;
  wire[46:0] T16975;
  wire[46:0] T16976;
  wire[44:0] T16977;
  wire[44:0] T16978;
  wire[1:0] T16979;
  wire T16980;
  wire T16981;
  wire T16982;
  wire[46:0] T16983;
  wire[46:0] T16984;
  wire[46:0] twiddle4_2_284_real;
  wire[46:0] T16985;
  wire[46:0] T16986;
  wire[46:0] T16987;
  wire[44:0] T16988;
  wire[44:0] T16989;
  wire[1:0] T16990;
  wire T16991;
  wire[46:0] twiddle4_2_285_real;
  wire[46:0] T16992;
  wire[46:0] T16993;
  wire[46:0] T16994;
  wire[44:0] T16995;
  wire[44:0] T16996;
  wire[1:0] T16997;
  wire T16998;
  wire T16999;
  wire[46:0] T17000;
  wire[46:0] twiddle4_2_286_real;
  wire[46:0] T17001;
  wire[46:0] T17002;
  wire[46:0] T17003;
  wire[44:0] T17004;
  wire[44:0] T17005;
  wire[1:0] T17006;
  wire T17007;
  wire[46:0] twiddle4_2_287_real;
  wire[46:0] T17008;
  wire[46:0] T17009;
  wire[46:0] T17010;
  wire[44:0] T17011;
  wire[44:0] T17012;
  wire[1:0] T17013;
  wire T17014;
  wire T17015;
  wire T17016;
  wire T17017;
  wire T17018;
  wire T17019;
  wire T17020;
  wire[47:0] T17021;
  wire[46:0] T17022;
  wire[46:0] T17023;
  wire[46:0] T17024;
  wire[46:0] T17025;
  wire[46:0] T17026;
  wire[46:0] twiddle4_2_288_real;
  wire[46:0] T17027;
  wire[46:0] T17028;
  wire[46:0] T17029;
  wire[44:0] T17030;
  wire[44:0] T17031;
  wire[1:0] T17032;
  wire T17033;
  wire[46:0] twiddle4_2_289_real;
  wire[46:0] T17034;
  wire[46:0] T17035;
  wire[46:0] T17036;
  wire[44:0] T17037;
  wire[44:0] T17038;
  wire[1:0] T17039;
  wire T17040;
  wire T17041;
  wire[46:0] T17042;
  wire[46:0] twiddle4_2_290_real;
  wire[46:0] T17043;
  wire[46:0] T17044;
  wire[46:0] T17045;
  wire[44:0] T17046;
  wire[44:0] T17047;
  wire[1:0] T17048;
  wire T17049;
  wire[46:0] twiddle4_2_291_real;
  wire[46:0] T17050;
  wire[46:0] T17051;
  wire[46:0] T17052;
  wire[44:0] T17053;
  wire[44:0] T17054;
  wire[1:0] T17055;
  wire T17056;
  wire T17057;
  wire T17058;
  wire[46:0] T17059;
  wire[46:0] T17060;
  wire[46:0] twiddle4_2_292_real;
  wire[46:0] T17061;
  wire[46:0] T17062;
  wire[46:0] T17063;
  wire[44:0] T17064;
  wire[44:0] T17065;
  wire[1:0] T17066;
  wire T17067;
  wire[46:0] twiddle4_2_293_real;
  wire[46:0] T17068;
  wire[46:0] T17069;
  wire[46:0] T17070;
  wire[44:0] T17071;
  wire[44:0] T17072;
  wire[1:0] T17073;
  wire T17074;
  wire T17075;
  wire[46:0] T17076;
  wire[46:0] twiddle4_2_294_real;
  wire[46:0] T17077;
  wire[46:0] T17078;
  wire[46:0] T17079;
  wire[44:0] T17080;
  wire[44:0] T17081;
  wire[1:0] T17082;
  wire T17083;
  wire[46:0] twiddle4_2_295_real;
  wire[46:0] T17084;
  wire[46:0] T17085;
  wire[46:0] T17086;
  wire[44:0] T17087;
  wire[44:0] T17088;
  wire[1:0] T17089;
  wire T17090;
  wire T17091;
  wire T17092;
  wire T17093;
  wire[46:0] T17094;
  wire[46:0] T17095;
  wire[46:0] T17096;
  wire[46:0] twiddle4_2_296_real;
  wire[46:0] T17097;
  wire[46:0] T17098;
  wire[46:0] T17099;
  wire[44:0] T17100;
  wire[44:0] T17101;
  wire[1:0] T17102;
  wire T17103;
  wire[46:0] twiddle4_2_297_real;
  wire[46:0] T17104;
  wire[46:0] T17105;
  wire[46:0] T17106;
  wire[44:0] T17107;
  wire[44:0] T17108;
  wire[1:0] T17109;
  wire T17110;
  wire T17111;
  wire[46:0] T17112;
  wire[46:0] twiddle4_2_298_real;
  wire[46:0] T17113;
  wire[46:0] T17114;
  wire[46:0] T17115;
  wire[45:0] T17116;
  wire[45:0] T17117;
  wire T17118;
  wire[46:0] twiddle4_2_299_real;
  wire[46:0] T17119;
  wire[46:0] T17120;
  wire[46:0] T17121;
  wire[45:0] T17122;
  wire[45:0] T17123;
  wire T17124;
  wire T17125;
  wire T17126;
  wire[46:0] T17127;
  wire[46:0] T17128;
  wire[46:0] twiddle4_2_300_real;
  wire[46:0] T17129;
  wire[46:0] T17130;
  wire[46:0] T17131;
  wire[45:0] T17132;
  wire[45:0] T17133;
  wire T17134;
  wire[46:0] twiddle4_2_301_real;
  wire[46:0] T17135;
  wire[46:0] T17136;
  wire[46:0] T17137;
  wire[45:0] T17138;
  wire[45:0] T17139;
  wire T17140;
  wire T17141;
  wire[46:0] T17142;
  wire[46:0] twiddle4_2_302_real;
  wire[46:0] T17143;
  wire[46:0] T17144;
  wire[46:0] T17145;
  wire[45:0] T17146;
  wire[45:0] T17147;
  wire T17148;
  wire[46:0] twiddle4_2_303_real;
  wire[46:0] T17149;
  wire[46:0] T17150;
  wire[46:0] T17151;
  wire[45:0] T17152;
  wire[45:0] T17153;
  wire T17154;
  wire T17155;
  wire T17156;
  wire T17157;
  wire T17158;
  wire[46:0] T17159;
  wire[46:0] T17160;
  wire[46:0] T17161;
  wire[46:0] T17162;
  wire[46:0] twiddle4_2_304_real;
  wire[46:0] T17163;
  wire[46:0] T17164;
  wire[46:0] T17165;
  wire[45:0] T17166;
  wire[45:0] T17167;
  wire T17168;
  wire[46:0] twiddle4_2_305_real;
  wire[46:0] T17169;
  wire[46:0] T17170;
  wire[46:0] T17171;
  wire[45:0] T17172;
  wire[45:0] T17173;
  wire T17174;
  wire T17175;
  wire[46:0] T17176;
  wire[46:0] twiddle4_2_306_real;
  wire[46:0] T17177;
  wire[46:0] T17178;
  wire[46:0] T17179;
  wire[45:0] T17180;
  wire[45:0] T17181;
  wire T17182;
  wire[46:0] twiddle4_2_307_real;
  wire[46:0] T17183;
  wire[46:0] T17184;
  wire[46:0] T17185;
  wire[45:0] T17186;
  wire[45:0] T17187;
  wire T17188;
  wire T17189;
  wire T17190;
  wire[46:0] T17191;
  wire[46:0] T17192;
  wire[46:0] twiddle4_2_308_real;
  wire[46:0] T17193;
  wire[46:0] T17194;
  wire[46:0] T17195;
  wire[45:0] T17196;
  wire[45:0] T17197;
  wire T17198;
  wire[46:0] twiddle4_2_309_real;
  wire[46:0] T17199;
  wire[46:0] T17200;
  wire[46:0] T17201;
  wire[45:0] T17202;
  wire[45:0] T17203;
  wire T17204;
  wire T17205;
  wire[46:0] T17206;
  wire[46:0] twiddle4_2_310_real;
  wire[46:0] T17207;
  wire[46:0] T17208;
  wire[46:0] T17209;
  wire[45:0] T17210;
  wire[45:0] T17211;
  wire T17212;
  wire[46:0] twiddle4_2_311_real;
  wire[46:0] T17213;
  wire[46:0] T17214;
  wire[46:0] T17215;
  wire[45:0] T17216;
  wire[45:0] T17217;
  wire T17218;
  wire T17219;
  wire T17220;
  wire T17221;
  wire[46:0] T17222;
  wire[46:0] T17223;
  wire[46:0] T17224;
  wire[46:0] twiddle4_2_312_real;
  wire[46:0] T17225;
  wire[46:0] T17226;
  wire[46:0] T17227;
  wire[45:0] T17228;
  wire[45:0] T17229;
  wire T17230;
  wire[46:0] twiddle4_2_313_real;
  wire[46:0] T17231;
  wire[46:0] T17232;
  wire[46:0] T17233;
  wire[45:0] T17234;
  wire[45:0] T17235;
  wire T17236;
  wire T17237;
  wire[46:0] T17238;
  wire[46:0] twiddle4_2_314_real;
  wire[46:0] T17239;
  wire[46:0] T17240;
  wire[46:0] T17241;
  wire[45:0] T17242;
  wire[45:0] T17243;
  wire T17244;
  wire[46:0] twiddle4_2_315_real;
  wire[46:0] T17245;
  wire[46:0] T17246;
  wire[46:0] T17247;
  wire[45:0] T17248;
  wire[45:0] T17249;
  wire T17250;
  wire T17251;
  wire T17252;
  wire[46:0] T17253;
  wire[46:0] T17254;
  wire[46:0] twiddle4_2_316_real;
  wire[46:0] T17255;
  wire[46:0] T17256;
  wire[46:0] T17257;
  wire[45:0] T17258;
  wire[45:0] T17259;
  wire T17260;
  wire[46:0] twiddle4_2_317_real;
  wire[46:0] T17261;
  wire[46:0] T17262;
  wire[46:0] T17263;
  wire[45:0] T17264;
  wire[45:0] T17265;
  wire T17266;
  wire T17267;
  wire[46:0] T17268;
  wire[46:0] twiddle4_2_318_real;
  wire[46:0] T17269;
  wire[46:0] T17270;
  wire[46:0] T17271;
  wire[45:0] T17272;
  wire[45:0] T17273;
  wire T17274;
  wire[46:0] twiddle4_2_319_real;
  wire[46:0] T17275;
  wire[46:0] T17276;
  wire[46:0] T17277;
  wire[45:0] T17278;
  wire[45:0] T17279;
  wire T17280;
  wire T17281;
  wire T17282;
  wire T17283;
  wire T17284;
  wire T17285;
  wire T17286;
  wire T17287;
  wire[47:0] T17288;
  wire[46:0] T17289;
  wire[46:0] T17290;
  wire[46:0] T17291;
  wire[46:0] T17292;
  wire[46:0] T17293;
  wire[46:0] T17294;
  wire[46:0] twiddle4_2_320_real;
  wire[46:0] T17295;
  wire[46:0] T17296;
  wire[46:0] T17297;
  wire[45:0] T17298;
  wire[45:0] T17299;
  wire T17300;
  wire[46:0] twiddle4_2_321_real;
  wire[46:0] T17301;
  wire[46:0] T17302;
  wire[46:0] T17303;
  wire[45:0] T17304;
  wire[45:0] T17305;
  wire T17306;
  wire T17307;
  wire[46:0] T17308;
  wire[46:0] twiddle4_2_322_real;
  wire[46:0] T17309;
  wire[46:0] T17310;
  wire[46:0] T17311;
  wire[45:0] T17312;
  wire[45:0] T17313;
  wire T17314;
  wire[46:0] twiddle4_2_323_real;
  wire[46:0] T17315;
  wire[46:0] T17316;
  wire[46:0] T17317;
  wire[45:0] T17318;
  wire[45:0] T17319;
  wire T17320;
  wire T17321;
  wire T17322;
  wire[46:0] T17323;
  wire[46:0] T17324;
  wire[46:0] twiddle4_2_324_real;
  wire[46:0] T17325;
  wire[46:0] T17326;
  wire[46:0] T17327;
  wire[45:0] T17328;
  wire[45:0] T17329;
  wire T17330;
  wire[46:0] twiddle4_2_325_real;
  wire[46:0] T17331;
  wire[46:0] T17332;
  wire[46:0] T17333;
  wire[45:0] T17334;
  wire[45:0] T17335;
  wire T17336;
  wire T17337;
  wire[46:0] T17338;
  wire[46:0] twiddle4_2_326_real;
  wire[46:0] T17339;
  wire[46:0] T17340;
  wire[46:0] T17341;
  wire[45:0] T17342;
  wire[45:0] T17343;
  wire T17344;
  wire[46:0] twiddle4_2_327_real;
  wire[46:0] T17345;
  wire[46:0] T17346;
  wire[46:0] T17347;
  wire[45:0] T17348;
  wire[45:0] T17349;
  wire T17350;
  wire T17351;
  wire T17352;
  wire T17353;
  wire[46:0] T17354;
  wire[46:0] T17355;
  wire[46:0] T17356;
  wire[46:0] twiddle4_2_328_real;
  wire[46:0] T17357;
  wire[46:0] T17358;
  wire[46:0] T17359;
  wire[45:0] T17360;
  wire[45:0] T17361;
  wire T17362;
  wire[46:0] twiddle4_2_329_real;
  wire[46:0] T17363;
  wire[46:0] T17364;
  wire[46:0] T17365;
  wire[45:0] T17366;
  wire[45:0] T17367;
  wire T17368;
  wire T17369;
  wire[46:0] T17370;
  wire[46:0] twiddle4_2_330_real;
  wire[46:0] T17371;
  wire[46:0] T17372;
  wire[46:0] T17373;
  wire[45:0] T17374;
  wire[45:0] T17375;
  wire T17376;
  wire[46:0] twiddle4_2_331_real;
  wire[46:0] T17377;
  wire[46:0] T17378;
  wire[46:0] T17379;
  wire[45:0] T17380;
  wire[45:0] T17381;
  wire T17382;
  wire T17383;
  wire T17384;
  wire[46:0] T17385;
  wire[46:0] T17386;
  wire[46:0] twiddle4_2_332_real;
  wire[46:0] T17387;
  wire[46:0] T17388;
  wire[46:0] T17389;
  wire[45:0] T17390;
  wire[45:0] T17391;
  wire T17392;
  wire[46:0] twiddle4_2_333_real;
  wire[46:0] T17393;
  wire[46:0] T17394;
  wire[46:0] T17395;
  wire[45:0] T17396;
  wire[45:0] T17397;
  wire T17398;
  wire T17399;
  wire[46:0] T17400;
  wire[46:0] twiddle4_2_334_real;
  wire[46:0] T17401;
  wire[46:0] T17402;
  wire[46:0] T17403;
  wire[45:0] T17404;
  wire[45:0] T17405;
  wire T17406;
  wire[46:0] twiddle4_2_335_real;
  wire[46:0] T17407;
  wire[46:0] T17408;
  wire[46:0] T17409;
  wire[45:0] T17410;
  wire[45:0] T17411;
  wire T17412;
  wire T17413;
  wire T17414;
  wire T17415;
  wire T17416;
  wire[46:0] T17417;
  wire[46:0] T17418;
  wire[46:0] T17419;
  wire[46:0] T17420;
  wire[46:0] twiddle4_2_336_real;
  wire[46:0] T17421;
  wire[46:0] T17422;
  wire[46:0] T17423;
  wire[45:0] T17424;
  wire[45:0] T17425;
  wire T17426;
  wire[46:0] twiddle4_2_337_real;
  wire[46:0] T17427;
  wire[46:0] T17428;
  wire[46:0] T17429;
  wire[45:0] T17430;
  wire[45:0] T17431;
  wire T17432;
  wire T17433;
  wire[46:0] T17434;
  wire[46:0] twiddle4_2_338_real;
  wire[46:0] T17435;
  wire[46:0] T17436;
  wire[46:0] T17437;
  wire[45:0] T17438;
  wire[45:0] T17439;
  wire T17440;
  wire[46:0] twiddle4_2_339_real;
  wire[46:0] T17441;
  wire[46:0] T17442;
  wire[46:0] T17443;
  wire[45:0] T17444;
  wire[45:0] T17445;
  wire T17446;
  wire T17447;
  wire T17448;
  wire[46:0] T17449;
  wire[46:0] T17450;
  wire[46:0] twiddle4_2_340_real;
  wire[46:0] T17451;
  wire[46:0] T17452;
  wire[46:0] T17453;
  wire[45:0] T17454;
  wire[45:0] T17455;
  wire T17456;
  wire[46:0] twiddle4_2_341_real;
  wire[46:0] T17457;
  wire[46:0] T17458;
  wire[46:0] T17459;
  wire[45:0] T17460;
  wire[45:0] T17461;
  wire T17462;
  wire T17463;
  wire[46:0] T17464;
  wire[46:0] twiddle4_2_342_real;
  wire[46:0] T17465;
  wire[46:0] T17466;
  wire[46:0] T17467;
  wire[46:0] T17468;
  wire[46:0] twiddle4_2_343_real;
  wire[46:0] T17469;
  wire[46:0] T17470;
  wire[46:0] T17471;
  wire[46:0] T17472;
  wire T17473;
  wire T17474;
  wire T17475;
  wire[46:0] T17476;
  wire[46:0] T17477;
  wire[46:0] T17478;
  wire[46:0] twiddle4_2_344_real;
  wire[46:0] T17479;
  wire[46:0] T17480;
  wire[46:0] T17481;
  wire[46:0] T17482;
  wire[46:0] twiddle4_2_345_real;
  wire[46:0] T17483;
  wire[46:0] T17484;
  wire[46:0] T17485;
  wire[46:0] T17486;
  wire T17487;
  wire[46:0] T17488;
  wire[46:0] twiddle4_2_346_real;
  wire[46:0] T17489;
  wire[46:0] T17490;
  wire[46:0] T17491;
  wire[46:0] T17492;
  wire[46:0] twiddle4_2_347_real;
  wire[46:0] T17493;
  wire[46:0] T17494;
  wire[46:0] T17495;
  wire[46:0] T17496;
  wire T17497;
  wire T17498;
  wire[46:0] T17499;
  wire[46:0] T17500;
  wire[46:0] twiddle4_2_348_real;
  wire[46:0] T17501;
  wire[46:0] T17502;
  wire[46:0] T17503;
  wire[46:0] T17504;
  wire[46:0] twiddle4_2_349_real;
  wire[46:0] T17505;
  wire[46:0] T17506;
  wire[46:0] T17507;
  wire[46:0] T17508;
  wire T17509;
  wire[46:0] T17510;
  wire[46:0] twiddle4_2_350_real;
  wire[46:0] T17511;
  wire[46:0] T17512;
  wire[46:0] T17513;
  wire[46:0] T17514;
  wire[46:0] twiddle4_2_351_real;
  wire[46:0] T17515;
  wire[46:0] T17516;
  wire[46:0] T17517;
  wire[46:0] T17518;
  wire T17519;
  wire T17520;
  wire T17521;
  wire T17522;
  wire T17523;
  wire[46:0] T17524;
  wire[46:0] T17525;
  wire[46:0] T17526;
  wire[46:0] T17527;
  wire[46:0] T17528;
  wire[46:0] twiddle4_2_352_real;
  wire[46:0] T17529;
  wire[46:0] T17530;
  wire[46:0] T17531;
  wire[46:0] T17532;
  wire[46:0] twiddle4_2_353_real;
  wire[46:0] T17533;
  wire[46:0] T17534;
  wire[46:0] T17535;
  wire[46:0] T17536;
  wire T17537;
  wire[46:0] T17538;
  wire[46:0] twiddle4_2_354_real;
  wire[46:0] T17539;
  wire[46:0] T17540;
  wire[46:0] T17541;
  wire[46:0] T17542;
  wire[46:0] twiddle4_2_355_real;
  wire[46:0] T17543;
  wire[46:0] T17544;
  wire[46:0] T17545;
  wire[46:0] T17546;
  wire T17547;
  wire T17548;
  wire[46:0] T17549;
  wire[46:0] T17550;
  wire[46:0] twiddle4_2_356_real;
  wire[46:0] T17551;
  wire[46:0] T17552;
  wire[46:0] T17553;
  wire[46:0] T17554;
  wire[46:0] twiddle4_2_357_real;
  wire[46:0] T17555;
  wire[46:0] T17556;
  wire[46:0] T17557;
  wire[46:0] T17558;
  wire T17559;
  wire[46:0] T17560;
  wire[46:0] twiddle4_2_358_real;
  wire[46:0] T17561;
  wire[46:0] T17562;
  wire[46:0] T17563;
  wire[46:0] T17564;
  wire[46:0] twiddle4_2_359_real;
  wire[46:0] T17565;
  wire[46:0] T17566;
  wire[46:0] T17567;
  wire[46:0] T17568;
  wire T17569;
  wire T17570;
  wire T17571;
  wire[46:0] T17572;
  wire[46:0] T17573;
  wire[46:0] T17574;
  wire[46:0] twiddle4_2_360_real;
  wire[46:0] T17575;
  wire[46:0] T17576;
  wire[46:0] T17577;
  wire[46:0] T17578;
  wire[46:0] twiddle4_2_361_real;
  wire[46:0] T17579;
  wire[46:0] T17580;
  wire[46:0] T17581;
  wire[46:0] T17582;
  wire T17583;
  wire[46:0] T17584;
  wire[46:0] twiddle4_2_362_real;
  wire[46:0] T17585;
  wire[46:0] T17586;
  wire[46:0] T17587;
  wire[46:0] T17588;
  wire[46:0] twiddle4_2_363_real;
  wire[46:0] T17589;
  wire[46:0] T17590;
  wire[46:0] T17591;
  wire[46:0] T17592;
  wire T17593;
  wire T17594;
  wire[46:0] T17595;
  wire[46:0] T17596;
  wire[46:0] twiddle4_2_364_real;
  wire[46:0] T17597;
  wire[46:0] T17598;
  wire[46:0] T17599;
  wire[46:0] T17600;
  wire[46:0] twiddle4_2_365_real;
  wire[46:0] T17601;
  wire[46:0] T17602;
  wire[46:0] T17603;
  wire[46:0] T17604;
  wire T17605;
  wire[46:0] T17606;
  wire[46:0] twiddle4_2_366_real;
  wire[46:0] T17607;
  wire[46:0] T17608;
  wire[46:0] T17609;
  wire[46:0] T17610;
  wire[46:0] twiddle4_2_367_real;
  wire[46:0] T17611;
  wire[46:0] T17612;
  wire[46:0] T17613;
  wire[46:0] T17614;
  wire T17615;
  wire T17616;
  wire T17617;
  wire T17618;
  wire[46:0] T17619;
  wire[46:0] T17620;
  wire[46:0] T17621;
  wire[46:0] T17622;
  wire[46:0] twiddle4_2_368_real;
  wire[46:0] T17623;
  wire[46:0] T17624;
  wire[46:0] T17625;
  wire[46:0] T17626;
  wire[46:0] twiddle4_2_369_real;
  wire[46:0] T17627;
  wire[46:0] T17628;
  wire[46:0] T17629;
  wire[46:0] T17630;
  wire T17631;
  wire[46:0] T17632;
  wire[46:0] twiddle4_2_370_real;
  wire[46:0] T17633;
  wire[46:0] T17634;
  wire[46:0] T17635;
  wire[46:0] T17636;
  wire[46:0] twiddle4_2_371_real;
  wire[46:0] T17637;
  wire[46:0] T17638;
  wire[46:0] T17639;
  wire[46:0] T17640;
  wire T17641;
  wire T17642;
  wire[46:0] T17643;
  wire[46:0] T17644;
  wire[46:0] twiddle4_2_372_real;
  wire[46:0] T17645;
  wire[46:0] T17646;
  wire[46:0] T17647;
  wire[46:0] T17648;
  wire[46:0] twiddle4_2_373_real;
  wire[46:0] T17649;
  wire[46:0] T17650;
  wire[46:0] T17651;
  wire[46:0] T17652;
  wire T17653;
  wire[46:0] T17654;
  wire[46:0] twiddle4_2_374_real;
  wire[46:0] T17655;
  wire[46:0] T17656;
  wire[46:0] T17657;
  wire[46:0] T17658;
  wire[46:0] twiddle4_2_375_real;
  wire[46:0] T17659;
  wire[46:0] T17660;
  wire[46:0] T17661;
  wire[46:0] T17662;
  wire T17663;
  wire T17664;
  wire T17665;
  wire[46:0] T17666;
  wire[46:0] T17667;
  wire[46:0] T17668;
  wire[46:0] twiddle4_2_376_real;
  wire[46:0] T17669;
  wire[46:0] T17670;
  wire[46:0] T17671;
  wire[46:0] T17672;
  wire[46:0] twiddle4_2_377_real;
  wire[46:0] T17673;
  wire[46:0] T17674;
  wire[46:0] T17675;
  wire[46:0] T17676;
  wire T17677;
  wire[46:0] T17678;
  wire[46:0] twiddle4_2_378_real;
  wire[46:0] T17679;
  wire[46:0] T17680;
  wire[46:0] T17681;
  wire[46:0] T17682;
  wire[46:0] twiddle4_2_379_real;
  wire[46:0] T17683;
  wire[46:0] T17684;
  wire[46:0] T17685;
  wire[46:0] T17686;
  wire T17687;
  wire T17688;
  wire[46:0] T17689;
  wire[46:0] T17690;
  wire[46:0] twiddle4_2_380_real;
  wire[46:0] T17691;
  wire[46:0] T17692;
  wire[46:0] T17693;
  wire[46:0] T17694;
  wire[46:0] twiddle4_2_381_real;
  wire[46:0] T17695;
  wire[46:0] T17696;
  wire[46:0] T17697;
  wire[46:0] T17698;
  wire T17699;
  wire[46:0] T17700;
  wire[46:0] twiddle4_2_382_real;
  wire[46:0] T17701;
  wire[46:0] T17702;
  wire[46:0] T17703;
  wire[46:0] T17704;
  wire[46:0] twiddle4_2_383_real;
  wire[46:0] T17705;
  wire[46:0] T17706;
  wire[46:0] T17707;
  wire[46:0] T17708;
  wire T17709;
  wire T17710;
  wire T17711;
  wire T17712;
  wire T17713;
  wire T17714;
  wire T17715;
  wire T17716;
  wire[47:0] T17717;
  wire[46:0] T17718;
  wire[46:0] T17719;
  wire[46:0] T17720;
  wire[46:0] T17721;
  wire[46:0] T17722;
  wire[46:0] T17723;
  wire[46:0] T17724;
  wire[46:0] twiddle4_2_384_real;
  wire[46:0] T17725;
  wire[46:0] T17726;
  wire[46:0] T17727;
  wire[46:0] T17728;
  wire[46:0] twiddle4_2_385_real;
  wire[46:0] T17729;
  wire[46:0] T17730;
  wire[46:0] T17731;
  wire[46:0] T17732;
  wire T17733;
  wire[46:0] T17734;
  wire[46:0] twiddle4_2_386_real;
  wire[46:0] T17735;
  wire[46:0] T17736;
  wire[46:0] T17737;
  wire[46:0] T17738;
  wire[46:0] twiddle4_2_387_real;
  wire[46:0] T17739;
  wire[46:0] T17740;
  wire[46:0] T17741;
  wire[46:0] T17742;
  wire T17743;
  wire T17744;
  wire[46:0] T17745;
  wire[46:0] T17746;
  wire[46:0] twiddle4_2_388_real;
  wire[46:0] T17747;
  wire[46:0] T17748;
  wire[46:0] T17749;
  wire[46:0] T17750;
  wire[46:0] twiddle4_2_389_real;
  wire[46:0] T17751;
  wire[46:0] T17752;
  wire[46:0] T17753;
  wire[46:0] T17754;
  wire T17755;
  wire[46:0] T17756;
  wire[46:0] twiddle4_2_390_real;
  wire[46:0] T17757;
  wire[46:0] T17758;
  wire[46:0] T17759;
  wire[46:0] T17760;
  wire[46:0] twiddle4_2_391_real;
  wire[46:0] T17761;
  wire[46:0] T17762;
  wire[46:0] T17763;
  wire[46:0] T17764;
  wire T17765;
  wire T17766;
  wire T17767;
  wire[46:0] T17768;
  wire[46:0] T17769;
  wire[46:0] T17770;
  wire[46:0] twiddle4_2_392_real;
  wire[46:0] T17771;
  wire[46:0] T17772;
  wire[46:0] T17773;
  wire[46:0] T17774;
  wire[46:0] twiddle4_2_393_real;
  wire[46:0] T17775;
  wire[46:0] T17776;
  wire[46:0] T17777;
  wire[46:0] T17778;
  wire T17779;
  wire[46:0] T17780;
  wire[46:0] twiddle4_2_394_real;
  wire[46:0] T17781;
  wire[46:0] T17782;
  wire[46:0] T17783;
  wire[46:0] T17784;
  wire[46:0] twiddle4_2_395_real;
  wire[46:0] T17785;
  wire[46:0] T17786;
  wire[46:0] T17787;
  wire[46:0] T17788;
  wire T17789;
  wire T17790;
  wire[46:0] T17791;
  wire[46:0] T17792;
  wire[46:0] twiddle4_2_396_real;
  wire[46:0] T17793;
  wire[46:0] T17794;
  wire[46:0] T17795;
  wire[46:0] T17796;
  wire[46:0] twiddle4_2_397_real;
  wire[46:0] T17797;
  wire[46:0] T17798;
  wire[46:0] T17799;
  wire[46:0] T17800;
  wire T17801;
  wire[46:0] T17802;
  wire[46:0] twiddle4_2_398_real;
  wire[46:0] T17803;
  wire[46:0] T17804;
  wire[46:0] T17805;
  wire[46:0] T17806;
  wire[46:0] twiddle4_2_399_real;
  wire[46:0] T17807;
  wire[46:0] T17808;
  wire[46:0] T17809;
  wire[46:0] T17810;
  wire T17811;
  wire T17812;
  wire T17813;
  wire T17814;
  wire[46:0] T17815;
  wire[46:0] T17816;
  wire[46:0] T17817;
  wire[46:0] T17818;
  wire[46:0] twiddle4_2_400_real;
  wire[46:0] T17819;
  wire[46:0] T17820;
  wire[46:0] T17821;
  wire[46:0] T17822;
  wire[46:0] twiddle4_2_401_real;
  wire[46:0] T17823;
  wire[46:0] T17824;
  wire[46:0] T17825;
  wire[46:0] T17826;
  wire T17827;
  wire[46:0] T17828;
  wire[46:0] twiddle4_2_402_real;
  wire[46:0] T17829;
  wire[46:0] T17830;
  wire[46:0] T17831;
  wire[46:0] T17832;
  wire[46:0] twiddle4_2_403_real;
  wire[46:0] T17833;
  wire[46:0] T17834;
  wire[46:0] T17835;
  wire[46:0] T17836;
  wire T17837;
  wire T17838;
  wire[46:0] T17839;
  wire[46:0] T17840;
  wire[46:0] twiddle4_2_404_real;
  wire[46:0] T17841;
  wire[46:0] T17842;
  wire[46:0] T17843;
  wire[46:0] T17844;
  wire[46:0] twiddle4_2_405_real;
  wire[46:0] T17845;
  wire[46:0] T17846;
  wire[46:0] T17847;
  wire[46:0] T17848;
  wire T17849;
  wire[46:0] T17850;
  wire[46:0] twiddle4_2_406_real;
  wire[46:0] T17851;
  wire[46:0] T17852;
  wire[46:0] T17853;
  wire[46:0] T17854;
  wire[46:0] twiddle4_2_407_real;
  wire[46:0] T17855;
  wire[46:0] T17856;
  wire[46:0] T17857;
  wire[46:0] T17858;
  wire T17859;
  wire T17860;
  wire T17861;
  wire[46:0] T17862;
  wire[46:0] T17863;
  wire[46:0] T17864;
  wire[46:0] twiddle4_2_408_real;
  wire[46:0] T17865;
  wire[46:0] T17866;
  wire[46:0] T17867;
  wire[46:0] T17868;
  wire[46:0] twiddle4_2_409_real;
  wire[46:0] T17869;
  wire[46:0] T17870;
  wire[46:0] T17871;
  wire[46:0] T17872;
  wire T17873;
  wire[46:0] T17874;
  wire[46:0] twiddle4_2_410_real;
  wire[46:0] T17875;
  wire[46:0] T17876;
  wire[46:0] T17877;
  wire[46:0] T17878;
  wire[46:0] twiddle4_2_411_real;
  wire[46:0] T17879;
  wire[46:0] T17880;
  wire[46:0] T17881;
  wire[46:0] T17882;
  wire T17883;
  wire T17884;
  wire[46:0] T17885;
  wire[46:0] T17886;
  wire[46:0] twiddle4_2_412_real;
  wire[46:0] T17887;
  wire[46:0] T17888;
  wire[46:0] T17889;
  wire[46:0] T17890;
  wire[46:0] twiddle4_2_413_real;
  wire[46:0] T17891;
  wire[46:0] T17892;
  wire[46:0] T17893;
  wire[46:0] T17894;
  wire T17895;
  wire[46:0] T17896;
  wire[46:0] twiddle4_2_414_real;
  wire[46:0] T17897;
  wire[46:0] T17898;
  wire[46:0] T17899;
  wire[46:0] T17900;
  wire[46:0] twiddle4_2_415_real;
  wire[46:0] T17901;
  wire[46:0] T17902;
  wire[46:0] T17903;
  wire[46:0] T17904;
  wire T17905;
  wire T17906;
  wire T17907;
  wire T17908;
  wire T17909;
  wire[46:0] T17910;
  wire[46:0] T17911;
  wire[46:0] T17912;
  wire[46:0] T17913;
  wire[46:0] T17914;
  wire[46:0] twiddle4_2_416_real;
  wire[46:0] T17915;
  wire[46:0] T17916;
  wire[46:0] T17917;
  wire[46:0] T17918;
  wire[46:0] twiddle4_2_417_real;
  wire[46:0] T17919;
  wire[46:0] T17920;
  wire[46:0] T17921;
  wire[46:0] T17922;
  wire T17923;
  wire[46:0] T17924;
  wire[46:0] twiddle4_2_418_real;
  wire[46:0] T17925;
  wire[46:0] T17926;
  wire[46:0] T17927;
  wire[46:0] T17928;
  wire[46:0] twiddle4_2_419_real;
  wire[46:0] T17929;
  wire[46:0] T17930;
  wire[46:0] T17931;
  wire[46:0] T17932;
  wire T17933;
  wire T17934;
  wire[46:0] T17935;
  wire[46:0] T17936;
  wire[46:0] twiddle4_2_420_real;
  wire[46:0] T17937;
  wire[46:0] T17938;
  wire[46:0] T17939;
  wire[46:0] T17940;
  wire[46:0] twiddle4_2_421_real;
  wire[46:0] T17941;
  wire[46:0] T17942;
  wire[46:0] T17943;
  wire[46:0] T17944;
  wire T17945;
  wire[46:0] T17946;
  wire[46:0] twiddle4_2_422_real;
  wire[46:0] T17947;
  wire[46:0] T17948;
  wire[46:0] T17949;
  wire[46:0] T17950;
  wire[46:0] twiddle4_2_423_real;
  wire[46:0] T17951;
  wire[46:0] T17952;
  wire[46:0] T17953;
  wire[46:0] T17954;
  wire T17955;
  wire T17956;
  wire T17957;
  wire[46:0] T17958;
  wire[46:0] T17959;
  wire[46:0] T17960;
  wire[46:0] twiddle4_2_424_real;
  wire[46:0] T17961;
  wire[46:0] T17962;
  wire[46:0] T17963;
  wire[46:0] T17964;
  wire[46:0] twiddle4_2_425_real;
  wire[46:0] T17965;
  wire[46:0] T17966;
  wire[46:0] T17967;
  wire[46:0] T17968;
  wire T17969;
  wire[46:0] T17970;
  wire[46:0] twiddle4_2_426_real;
  wire[46:0] T17971;
  wire[46:0] T17972;
  wire[46:0] T17973;
  wire[46:0] T17974;
  wire[46:0] twiddle4_2_427_real;
  wire[46:0] T17975;
  wire[45:0] T17976;
  wire[45:0] T17977;
  wire T17978;
  wire[46:0] T17979;
  wire[46:0] T17980;
  wire T17981;
  wire T17982;
  wire[46:0] T17983;
  wire[46:0] T17984;
  wire[46:0] twiddle4_2_428_real;
  wire[46:0] T17985;
  wire[45:0] T17986;
  wire[45:0] T17987;
  wire T17988;
  wire[46:0] T17989;
  wire[46:0] T17990;
  wire[46:0] twiddle4_2_429_real;
  wire[46:0] T17991;
  wire[45:0] T17992;
  wire[45:0] T17993;
  wire T17994;
  wire[46:0] T17995;
  wire[46:0] T17996;
  wire T17997;
  wire[46:0] T17998;
  wire[46:0] twiddle4_2_430_real;
  wire[46:0] T17999;
  wire[45:0] T18000;
  wire[45:0] T18001;
  wire T18002;
  wire[46:0] T18003;
  wire[46:0] T18004;
  wire[46:0] twiddle4_2_431_real;
  wire[46:0] T18005;
  wire[45:0] T18006;
  wire[45:0] T18007;
  wire T18008;
  wire[46:0] T18009;
  wire[46:0] T18010;
  wire T18011;
  wire T18012;
  wire T18013;
  wire T18014;
  wire[46:0] T18015;
  wire[46:0] T18016;
  wire[46:0] T18017;
  wire[46:0] T18018;
  wire[46:0] twiddle4_2_432_real;
  wire[46:0] T18019;
  wire[45:0] T18020;
  wire[45:0] T18021;
  wire T18022;
  wire[46:0] T18023;
  wire[46:0] T18024;
  wire[46:0] twiddle4_2_433_real;
  wire[46:0] T18025;
  wire[45:0] T18026;
  wire[45:0] T18027;
  wire T18028;
  wire[46:0] T18029;
  wire[46:0] T18030;
  wire T18031;
  wire[46:0] T18032;
  wire[46:0] twiddle4_2_434_real;
  wire[46:0] T18033;
  wire[45:0] T18034;
  wire[45:0] T18035;
  wire T18036;
  wire[46:0] T18037;
  wire[46:0] T18038;
  wire[46:0] twiddle4_2_435_real;
  wire[46:0] T18039;
  wire[45:0] T18040;
  wire[45:0] T18041;
  wire T18042;
  wire[46:0] T18043;
  wire[46:0] T18044;
  wire T18045;
  wire T18046;
  wire[46:0] T18047;
  wire[46:0] T18048;
  wire[46:0] twiddle4_2_436_real;
  wire[46:0] T18049;
  wire[45:0] T18050;
  wire[45:0] T18051;
  wire T18052;
  wire[46:0] T18053;
  wire[46:0] T18054;
  wire[46:0] twiddle4_2_437_real;
  wire[46:0] T18055;
  wire[45:0] T18056;
  wire[45:0] T18057;
  wire T18058;
  wire[46:0] T18059;
  wire[46:0] T18060;
  wire T18061;
  wire[46:0] T18062;
  wire[46:0] twiddle4_2_438_real;
  wire[46:0] T18063;
  wire[45:0] T18064;
  wire[45:0] T18065;
  wire T18066;
  wire[46:0] T18067;
  wire[46:0] T18068;
  wire[46:0] twiddle4_2_439_real;
  wire[46:0] T18069;
  wire[45:0] T18070;
  wire[45:0] T18071;
  wire T18072;
  wire[46:0] T18073;
  wire[46:0] T18074;
  wire T18075;
  wire T18076;
  wire T18077;
  wire[46:0] T18078;
  wire[46:0] T18079;
  wire[46:0] T18080;
  wire[46:0] twiddle4_2_440_real;
  wire[46:0] T18081;
  wire[45:0] T18082;
  wire[45:0] T18083;
  wire T18084;
  wire[46:0] T18085;
  wire[46:0] T18086;
  wire[46:0] twiddle4_2_441_real;
  wire[46:0] T18087;
  wire[45:0] T18088;
  wire[45:0] T18089;
  wire T18090;
  wire[46:0] T18091;
  wire[46:0] T18092;
  wire T18093;
  wire[46:0] T18094;
  wire[46:0] twiddle4_2_442_real;
  wire[46:0] T18095;
  wire[45:0] T18096;
  wire[45:0] T18097;
  wire T18098;
  wire[46:0] T18099;
  wire[46:0] T18100;
  wire[46:0] twiddle4_2_443_real;
  wire[46:0] T18101;
  wire[45:0] T18102;
  wire[45:0] T18103;
  wire T18104;
  wire[46:0] T18105;
  wire[46:0] T18106;
  wire T18107;
  wire T18108;
  wire[46:0] T18109;
  wire[46:0] T18110;
  wire[46:0] twiddle4_2_444_real;
  wire[46:0] T18111;
  wire[45:0] T18112;
  wire[45:0] T18113;
  wire T18114;
  wire[46:0] T18115;
  wire[46:0] T18116;
  wire[46:0] twiddle4_2_445_real;
  wire[46:0] T18117;
  wire[45:0] T18118;
  wire[45:0] T18119;
  wire T18120;
  wire[46:0] T18121;
  wire[46:0] T18122;
  wire T18123;
  wire[46:0] T18124;
  wire[46:0] twiddle4_2_446_real;
  wire[46:0] T18125;
  wire[45:0] T18126;
  wire[45:0] T18127;
  wire T18128;
  wire[46:0] T18129;
  wire[46:0] T18130;
  wire[46:0] twiddle4_2_447_real;
  wire[46:0] T18131;
  wire[45:0] T18132;
  wire[45:0] T18133;
  wire T18134;
  wire[46:0] T18135;
  wire[46:0] T18136;
  wire T18137;
  wire T18138;
  wire T18139;
  wire T18140;
  wire T18141;
  wire T18142;
  wire[46:0] T18143;
  wire[46:0] T18144;
  wire[46:0] T18145;
  wire[46:0] T18146;
  wire[46:0] T18147;
  wire[46:0] T18148;
  wire[46:0] twiddle4_2_448_real;
  wire[46:0] T18149;
  wire[45:0] T18150;
  wire[45:0] T18151;
  wire T18152;
  wire[46:0] T18153;
  wire[46:0] T18154;
  wire[46:0] twiddle4_2_449_real;
  wire[46:0] T18155;
  wire[45:0] T18156;
  wire[45:0] T18157;
  wire T18158;
  wire[46:0] T18159;
  wire[46:0] T18160;
  wire T18161;
  wire[46:0] T18162;
  wire[46:0] twiddle4_2_450_real;
  wire[46:0] T18163;
  wire[45:0] T18164;
  wire[45:0] T18165;
  wire T18166;
  wire[46:0] T18167;
  wire[46:0] T18168;
  wire[46:0] twiddle4_2_451_real;
  wire[46:0] T18169;
  wire[45:0] T18170;
  wire[45:0] T18171;
  wire T18172;
  wire[46:0] T18173;
  wire[46:0] T18174;
  wire T18175;
  wire T18176;
  wire[46:0] T18177;
  wire[46:0] T18178;
  wire[46:0] twiddle4_2_452_real;
  wire[46:0] T18179;
  wire[45:0] T18180;
  wire[45:0] T18181;
  wire T18182;
  wire[46:0] T18183;
  wire[46:0] T18184;
  wire[46:0] twiddle4_2_453_real;
  wire[46:0] T18185;
  wire[45:0] T18186;
  wire[45:0] T18187;
  wire T18188;
  wire[46:0] T18189;
  wire[46:0] T18190;
  wire T18191;
  wire[46:0] T18192;
  wire[46:0] twiddle4_2_454_real;
  wire[46:0] T18193;
  wire[45:0] T18194;
  wire[45:0] T18195;
  wire T18196;
  wire[46:0] T18197;
  wire[46:0] T18198;
  wire[46:0] twiddle4_2_455_real;
  wire[46:0] T18199;
  wire[45:0] T18200;
  wire[45:0] T18201;
  wire T18202;
  wire[46:0] T18203;
  wire[46:0] T18204;
  wire T18205;
  wire T18206;
  wire T18207;
  wire[46:0] T18208;
  wire[46:0] T18209;
  wire[46:0] T18210;
  wire[46:0] twiddle4_2_456_real;
  wire[46:0] T18211;
  wire[45:0] T18212;
  wire[45:0] T18213;
  wire T18214;
  wire[46:0] T18215;
  wire[46:0] T18216;
  wire[46:0] twiddle4_2_457_real;
  wire[46:0] T18217;
  wire[45:0] T18218;
  wire[45:0] T18219;
  wire T18220;
  wire[46:0] T18221;
  wire[46:0] T18222;
  wire T18223;
  wire[46:0] T18224;
  wire[46:0] twiddle4_2_458_real;
  wire[46:0] T18225;
  wire[45:0] T18226;
  wire[45:0] T18227;
  wire T18228;
  wire[46:0] T18229;
  wire[46:0] T18230;
  wire[46:0] twiddle4_2_459_real;
  wire[46:0] T18231;
  wire[45:0] T18232;
  wire[45:0] T18233;
  wire T18234;
  wire[46:0] T18235;
  wire[46:0] T18236;
  wire T18237;
  wire T18238;
  wire[46:0] T18239;
  wire[46:0] T18240;
  wire[46:0] twiddle4_2_460_real;
  wire[46:0] T18241;
  wire[45:0] T18242;
  wire[45:0] T18243;
  wire T18244;
  wire[46:0] T18245;
  wire[46:0] T18246;
  wire[46:0] twiddle4_2_461_real;
  wire[46:0] T18247;
  wire[45:0] T18248;
  wire[45:0] T18249;
  wire T18250;
  wire[46:0] T18251;
  wire[46:0] T18252;
  wire T18253;
  wire[46:0] T18254;
  wire[46:0] twiddle4_2_462_real;
  wire[46:0] T18255;
  wire[45:0] T18256;
  wire[45:0] T18257;
  wire T18258;
  wire[46:0] T18259;
  wire[46:0] T18260;
  wire[46:0] twiddle4_2_463_real;
  wire[46:0] T18261;
  wire[45:0] T18262;
  wire[45:0] T18263;
  wire T18264;
  wire[46:0] T18265;
  wire[46:0] T18266;
  wire T18267;
  wire T18268;
  wire T18269;
  wire T18270;
  wire[46:0] T18271;
  wire[46:0] T18272;
  wire[46:0] T18273;
  wire[46:0] T18274;
  wire[46:0] twiddle4_2_464_real;
  wire[46:0] T18275;
  wire[45:0] T18276;
  wire[45:0] T18277;
  wire T18278;
  wire[46:0] T18279;
  wire[46:0] T18280;
  wire[46:0] twiddle4_2_465_real;
  wire[46:0] T18281;
  wire[45:0] T18282;
  wire[45:0] T18283;
  wire T18284;
  wire[46:0] T18285;
  wire[46:0] T18286;
  wire T18287;
  wire[46:0] T18288;
  wire[46:0] twiddle4_2_466_real;
  wire[46:0] T18289;
  wire[45:0] T18290;
  wire[45:0] T18291;
  wire T18292;
  wire[46:0] T18293;
  wire[46:0] T18294;
  wire[46:0] twiddle4_2_467_real;
  wire[46:0] T18295;
  wire[45:0] T18296;
  wire[45:0] T18297;
  wire T18298;
  wire[46:0] T18299;
  wire[46:0] T18300;
  wire T18301;
  wire T18302;
  wire[46:0] T18303;
  wire[46:0] T18304;
  wire[46:0] twiddle4_2_468_real;
  wire[46:0] T18305;
  wire[45:0] T18306;
  wire[45:0] T18307;
  wire T18308;
  wire[46:0] T18309;
  wire[46:0] T18310;
  wire[46:0] twiddle4_2_469_real;
  wire[46:0] T18311;
  wire[45:0] T18312;
  wire[45:0] T18313;
  wire T18314;
  wire[46:0] T18315;
  wire[46:0] T18316;
  wire T18317;
  wire[46:0] T18318;
  wire[46:0] twiddle4_2_470_real;
  wire[46:0] T18319;
  wire[45:0] T18320;
  wire[45:0] T18321;
  wire T18322;
  wire[46:0] T18323;
  wire[46:0] T18324;
  wire[46:0] twiddle4_2_471_real;
  wire[46:0] T18325;
  wire[44:0] T18326;
  wire[44:0] T18327;
  wire[1:0] T18328;
  wire T18329;
  wire[46:0] T18330;
  wire[46:0] T18331;
  wire T18332;
  wire T18333;
  wire T18334;
  wire[46:0] T18335;
  wire[46:0] T18336;
  wire[46:0] T18337;
  wire[46:0] twiddle4_2_472_real;
  wire[46:0] T18338;
  wire[44:0] T18339;
  wire[44:0] T18340;
  wire[1:0] T18341;
  wire T18342;
  wire[46:0] T18343;
  wire[46:0] T18344;
  wire[46:0] twiddle4_2_473_real;
  wire[46:0] T18345;
  wire[44:0] T18346;
  wire[44:0] T18347;
  wire[1:0] T18348;
  wire T18349;
  wire[46:0] T18350;
  wire[46:0] T18351;
  wire T18352;
  wire[46:0] T18353;
  wire[46:0] twiddle4_2_474_real;
  wire[46:0] T18354;
  wire[44:0] T18355;
  wire[44:0] T18356;
  wire[1:0] T18357;
  wire T18358;
  wire[46:0] T18359;
  wire[46:0] T18360;
  wire[46:0] twiddle4_2_475_real;
  wire[46:0] T18361;
  wire[44:0] T18362;
  wire[44:0] T18363;
  wire[1:0] T18364;
  wire T18365;
  wire[46:0] T18366;
  wire[46:0] T18367;
  wire T18368;
  wire T18369;
  wire[46:0] T18370;
  wire[46:0] T18371;
  wire[46:0] twiddle4_2_476_real;
  wire[46:0] T18372;
  wire[44:0] T18373;
  wire[44:0] T18374;
  wire[1:0] T18375;
  wire T18376;
  wire[46:0] T18377;
  wire[46:0] T18378;
  wire[46:0] twiddle4_2_477_real;
  wire[46:0] T18379;
  wire[44:0] T18380;
  wire[44:0] T18381;
  wire[1:0] T18382;
  wire T18383;
  wire[46:0] T18384;
  wire[46:0] T18385;
  wire T18386;
  wire[46:0] T18387;
  wire[46:0] twiddle4_2_478_real;
  wire[46:0] T18388;
  wire[44:0] T18389;
  wire[44:0] T18390;
  wire[1:0] T18391;
  wire T18392;
  wire[46:0] T18393;
  wire[46:0] T18394;
  wire[46:0] twiddle4_2_479_real;
  wire[46:0] T18395;
  wire[44:0] T18396;
  wire[44:0] T18397;
  wire[1:0] T18398;
  wire T18399;
  wire[46:0] T18400;
  wire[46:0] T18401;
  wire T18402;
  wire T18403;
  wire T18404;
  wire T18405;
  wire T18406;
  wire[46:0] T18407;
  wire[46:0] T18408;
  wire[46:0] T18409;
  wire[46:0] T18410;
  wire[46:0] T18411;
  wire[46:0] twiddle4_2_480_real;
  wire[46:0] T18412;
  wire[44:0] T18413;
  wire[44:0] T18414;
  wire[1:0] T18415;
  wire T18416;
  wire[46:0] T18417;
  wire[46:0] T18418;
  wire[46:0] twiddle4_2_481_real;
  wire[46:0] T18419;
  wire[44:0] T18420;
  wire[44:0] T18421;
  wire[1:0] T18422;
  wire T18423;
  wire[46:0] T18424;
  wire[46:0] T18425;
  wire T18426;
  wire[46:0] T18427;
  wire[46:0] twiddle4_2_482_real;
  wire[46:0] T18428;
  wire[44:0] T18429;
  wire[44:0] T18430;
  wire[1:0] T18431;
  wire T18432;
  wire[46:0] T18433;
  wire[46:0] T18434;
  wire[46:0] twiddle4_2_483_real;
  wire[46:0] T18435;
  wire[44:0] T18436;
  wire[44:0] T18437;
  wire[1:0] T18438;
  wire T18439;
  wire[46:0] T18440;
  wire[46:0] T18441;
  wire T18442;
  wire T18443;
  wire[46:0] T18444;
  wire[46:0] T18445;
  wire[46:0] twiddle4_2_484_real;
  wire[46:0] T18446;
  wire[44:0] T18447;
  wire[44:0] T18448;
  wire[1:0] T18449;
  wire T18450;
  wire[46:0] T18451;
  wire[46:0] T18452;
  wire[46:0] twiddle4_2_485_real;
  wire[46:0] T18453;
  wire[44:0] T18454;
  wire[44:0] T18455;
  wire[1:0] T18456;
  wire T18457;
  wire[46:0] T18458;
  wire[46:0] T18459;
  wire T18460;
  wire[46:0] T18461;
  wire[46:0] twiddle4_2_486_real;
  wire[46:0] T18462;
  wire[44:0] T18463;
  wire[44:0] T18464;
  wire[1:0] T18465;
  wire T18466;
  wire[46:0] T18467;
  wire[46:0] T18468;
  wire[46:0] twiddle4_2_487_real;
  wire[46:0] T18469;
  wire[44:0] T18470;
  wire[44:0] T18471;
  wire[1:0] T18472;
  wire T18473;
  wire[46:0] T18474;
  wire[46:0] T18475;
  wire T18476;
  wire T18477;
  wire T18478;
  wire[46:0] T18479;
  wire[46:0] T18480;
  wire[46:0] T18481;
  wire[46:0] twiddle4_2_488_real;
  wire[46:0] T18482;
  wire[44:0] T18483;
  wire[44:0] T18484;
  wire[1:0] T18485;
  wire T18486;
  wire[46:0] T18487;
  wire[46:0] T18488;
  wire[46:0] twiddle4_2_489_real;
  wire[46:0] T18489;
  wire[44:0] T18490;
  wire[44:0] T18491;
  wire[1:0] T18492;
  wire T18493;
  wire[46:0] T18494;
  wire[46:0] T18495;
  wire T18496;
  wire[46:0] T18497;
  wire[46:0] twiddle4_2_490_real;
  wire[46:0] T18498;
  wire[44:0] T18499;
  wire[44:0] T18500;
  wire[1:0] T18501;
  wire T18502;
  wire[46:0] T18503;
  wire[46:0] T18504;
  wire[46:0] twiddle4_2_491_real;
  wire[46:0] T18505;
  wire[44:0] T18506;
  wire[44:0] T18507;
  wire[1:0] T18508;
  wire T18509;
  wire[46:0] T18510;
  wire[46:0] T18511;
  wire T18512;
  wire T18513;
  wire[46:0] T18514;
  wire[46:0] T18515;
  wire[46:0] twiddle4_2_492_real;
  wire[46:0] T18516;
  wire[43:0] T18517;
  wire[43:0] T18518;
  wire[2:0] T18519;
  wire T18520;
  wire[46:0] T18521;
  wire[46:0] T18522;
  wire[46:0] twiddle4_2_493_real;
  wire[46:0] T18523;
  wire[43:0] T18524;
  wire[43:0] T18525;
  wire[2:0] T18526;
  wire T18527;
  wire[46:0] T18528;
  wire[46:0] T18529;
  wire T18530;
  wire[46:0] T18531;
  wire[46:0] twiddle4_2_494_real;
  wire[46:0] T18532;
  wire[43:0] T18533;
  wire[43:0] T18534;
  wire[2:0] T18535;
  wire T18536;
  wire[46:0] T18537;
  wire[46:0] T18538;
  wire[46:0] twiddle4_2_495_real;
  wire[46:0] T18539;
  wire[43:0] T18540;
  wire[43:0] T18541;
  wire[2:0] T18542;
  wire T18543;
  wire[46:0] T18544;
  wire[46:0] T18545;
  wire T18546;
  wire T18547;
  wire T18548;
  wire T18549;
  wire[46:0] T18550;
  wire[46:0] T18551;
  wire[46:0] T18552;
  wire[46:0] T18553;
  wire[46:0] twiddle4_2_496_real;
  wire[46:0] T18554;
  wire[43:0] T18555;
  wire[43:0] T18556;
  wire[2:0] T18557;
  wire T18558;
  wire[46:0] T18559;
  wire[46:0] T18560;
  wire[46:0] twiddle4_2_497_real;
  wire[46:0] T18561;
  wire[43:0] T18562;
  wire[43:0] T18563;
  wire[2:0] T18564;
  wire T18565;
  wire[46:0] T18566;
  wire[46:0] T18567;
  wire T18568;
  wire[46:0] T18569;
  wire[46:0] twiddle4_2_498_real;
  wire[46:0] T18570;
  wire[43:0] T18571;
  wire[43:0] T18572;
  wire[2:0] T18573;
  wire T18574;
  wire[46:0] T18575;
  wire[46:0] T18576;
  wire[46:0] twiddle4_2_499_real;
  wire[46:0] T18577;
  wire[43:0] T18578;
  wire[43:0] T18579;
  wire[2:0] T18580;
  wire T18581;
  wire[46:0] T18582;
  wire[46:0] T18583;
  wire T18584;
  wire T18585;
  wire[46:0] T18586;
  wire[46:0] T18587;
  wire[46:0] twiddle4_2_500_real;
  wire[46:0] T18588;
  wire[43:0] T18589;
  wire[43:0] T18590;
  wire[2:0] T18591;
  wire T18592;
  wire[46:0] T18593;
  wire[46:0] T18594;
  wire[46:0] twiddle4_2_501_real;
  wire[46:0] T18595;
  wire[43:0] T18596;
  wire[43:0] T18597;
  wire[2:0] T18598;
  wire T18599;
  wire[46:0] T18600;
  wire[46:0] T18601;
  wire T18602;
  wire[46:0] T18603;
  wire[46:0] twiddle4_2_502_real;
  wire[46:0] T18604;
  wire[42:0] T18605;
  wire[42:0] T18606;
  wire[3:0] T18607;
  wire T18608;
  wire[46:0] T18609;
  wire[46:0] T18610;
  wire[46:0] twiddle4_2_503_real;
  wire[46:0] T18611;
  wire[42:0] T18612;
  wire[42:0] T18613;
  wire[3:0] T18614;
  wire T18615;
  wire[46:0] T18616;
  wire[46:0] T18617;
  wire T18618;
  wire T18619;
  wire T18620;
  wire[46:0] T18621;
  wire[46:0] T18622;
  wire[46:0] T18623;
  wire[46:0] twiddle4_2_504_real;
  wire[46:0] T18624;
  wire[42:0] T18625;
  wire[42:0] T18626;
  wire[3:0] T18627;
  wire T18628;
  wire[46:0] T18629;
  wire[46:0] T18630;
  wire[46:0] twiddle4_2_505_real;
  wire[46:0] T18631;
  wire[42:0] T18632;
  wire[42:0] T18633;
  wire[3:0] T18634;
  wire T18635;
  wire[46:0] T18636;
  wire[46:0] T18637;
  wire T18638;
  wire[46:0] T18639;
  wire[46:0] twiddle4_2_506_real;
  wire[46:0] T18640;
  wire[42:0] T18641;
  wire[42:0] T18642;
  wire[3:0] T18643;
  wire T18644;
  wire[46:0] T18645;
  wire[46:0] T18646;
  wire[46:0] twiddle4_2_507_real;
  wire[46:0] T18647;
  wire[41:0] T18648;
  wire[41:0] T18649;
  wire[4:0] T18650;
  wire T18651;
  wire[46:0] T18652;
  wire[46:0] T18653;
  wire T18654;
  wire T18655;
  wire[46:0] T18656;
  wire[46:0] T18657;
  wire[46:0] twiddle4_2_508_real;
  wire[46:0] T18658;
  wire[41:0] T18659;
  wire[41:0] T18660;
  wire[4:0] T18661;
  wire T18662;
  wire[46:0] T18663;
  wire[46:0] T18664;
  wire[46:0] twiddle4_2_509_real;
  wire[46:0] T18665;
  wire[41:0] T18666;
  wire[41:0] T18667;
  wire[4:0] T18668;
  wire T18669;
  wire[46:0] T18670;
  wire[46:0] T18671;
  wire T18672;
  wire[46:0] T18673;
  wire[46:0] twiddle4_2_510_real;
  wire[46:0] T18674;
  wire[40:0] T18675;
  wire[40:0] T18676;
  wire[5:0] T18677;
  wire T18678;
  wire[46:0] T18679;
  wire[46:0] T18680;
  wire[46:0] twiddle4_2_511_real;
  wire[46:0] T18681;
  wire[39:0] T18682;
  wire[39:0] T18683;
  wire[6:0] T18684;
  wire T18685;
  wire[46:0] T18686;
  wire[46:0] T18687;
  wire T18688;
  wire T18689;
  wire T18690;
  wire T18691;
  wire T18692;
  wire T18693;
  wire T18694;
  wire T18695;
  wire T18696;
  wire T18697;
  wire[15:0] T18698;
  wire[47:0] T18699;
  wire[47:0] T18700;
  wire[47:0] T18701;
  wire[47:0] T18702;
  wire[47:0] T18703;
  wire[47:0] T18704;
  wire[47:0] T18705;
  wire[47:0] T18706;
  wire[47:0] T18707;
  wire[47:0] twiddle4_1_0_imag;
  wire[47:0] T18708;
  wire[16:0] T18709;
  wire[16:0] T18710;
  wire[30:0] T18711;
  wire T18712;
  wire[47:0] T18713;
  wire[47:0] T18714;
  wire[47:0] T18715;
  wire[46:0] twiddle4_1_1_imag;
  wire[46:0] T18716;
  wire[38:0] T18717;
  wire[38:0] T18718;
  wire[7:0] T18719;
  wire T18720;
  wire[46:0] T18721;
  wire[46:0] T18722;
  wire T18723;
  wire T18724;
  wire[8:0] T18725;
  wire[8:0] T18726;
  wire[47:0] T18727;
  wire[46:0] T18728;
  wire[46:0] twiddle4_1_2_imag;
  wire[46:0] T18729;
  wire[39:0] T18730;
  wire[39:0] T18731;
  wire[6:0] T18732;
  wire T18733;
  wire[46:0] T18734;
  wire[46:0] T18735;
  wire[46:0] twiddle4_1_3_imag;
  wire[46:0] T18736;
  wire[40:0] T18737;
  wire[40:0] T18738;
  wire[5:0] T18739;
  wire T18740;
  wire[46:0] T18741;
  wire[46:0] T18742;
  wire T18743;
  wire T18744;
  wire T18745;
  wire[47:0] T18746;
  wire[46:0] T18747;
  wire[46:0] T18748;
  wire[46:0] twiddle4_1_4_imag;
  wire[46:0] T18749;
  wire[40:0] T18750;
  wire[40:0] T18751;
  wire[5:0] T18752;
  wire T18753;
  wire[46:0] T18754;
  wire[46:0] T18755;
  wire[46:0] twiddle4_1_5_imag;
  wire[46:0] T18756;
  wire[40:0] T18757;
  wire[40:0] T18758;
  wire[5:0] T18759;
  wire T18760;
  wire[46:0] T18761;
  wire[46:0] T18762;
  wire T18763;
  wire[46:0] T18764;
  wire[46:0] twiddle4_1_6_imag;
  wire[46:0] T18765;
  wire[41:0] T18766;
  wire[41:0] T18767;
  wire[4:0] T18768;
  wire T18769;
  wire[46:0] T18770;
  wire[46:0] T18771;
  wire[46:0] twiddle4_1_7_imag;
  wire[46:0] T18772;
  wire[41:0] T18773;
  wire[41:0] T18774;
  wire[4:0] T18775;
  wire T18776;
  wire[46:0] T18777;
  wire[46:0] T18778;
  wire T18779;
  wire T18780;
  wire T18781;
  wire T18782;
  wire[47:0] T18783;
  wire[46:0] T18784;
  wire[46:0] T18785;
  wire[46:0] T18786;
  wire[46:0] twiddle4_1_8_imag;
  wire[46:0] T18787;
  wire[41:0] T18788;
  wire[41:0] T18789;
  wire[4:0] T18790;
  wire T18791;
  wire[46:0] T18792;
  wire[46:0] T18793;
  wire[46:0] twiddle4_1_9_imag;
  wire[46:0] T18794;
  wire[41:0] T18795;
  wire[41:0] T18796;
  wire[4:0] T18797;
  wire T18798;
  wire[46:0] T18799;
  wire[46:0] T18800;
  wire T18801;
  wire[46:0] T18802;
  wire[46:0] twiddle4_1_10_imag;
  wire[46:0] T18803;
  wire[41:0] T18804;
  wire[41:0] T18805;
  wire[4:0] T18806;
  wire T18807;
  wire[46:0] T18808;
  wire[46:0] T18809;
  wire[46:0] twiddle4_1_11_imag;
  wire[46:0] T18810;
  wire[42:0] T18811;
  wire[42:0] T18812;
  wire[3:0] T18813;
  wire T18814;
  wire[46:0] T18815;
  wire[46:0] T18816;
  wire T18817;
  wire T18818;
  wire[46:0] T18819;
  wire[46:0] T18820;
  wire[46:0] twiddle4_1_12_imag;
  wire[46:0] T18821;
  wire[42:0] T18822;
  wire[42:0] T18823;
  wire[3:0] T18824;
  wire T18825;
  wire[46:0] T18826;
  wire[46:0] T18827;
  wire[46:0] twiddle4_1_13_imag;
  wire[46:0] T18828;
  wire[42:0] T18829;
  wire[42:0] T18830;
  wire[3:0] T18831;
  wire T18832;
  wire[46:0] T18833;
  wire[46:0] T18834;
  wire T18835;
  wire[46:0] T18836;
  wire[46:0] twiddle4_1_14_imag;
  wire[46:0] T18837;
  wire[42:0] T18838;
  wire[42:0] T18839;
  wire[3:0] T18840;
  wire T18841;
  wire[46:0] T18842;
  wire[46:0] T18843;
  wire[46:0] twiddle4_1_15_imag;
  wire[46:0] T18844;
  wire[42:0] T18845;
  wire[42:0] T18846;
  wire[3:0] T18847;
  wire T18848;
  wire[46:0] T18849;
  wire[46:0] T18850;
  wire T18851;
  wire T18852;
  wire T18853;
  wire T18854;
  wire T18855;
  wire[47:0] T18856;
  wire[46:0] T18857;
  wire[46:0] T18858;
  wire[46:0] T18859;
  wire[46:0] T18860;
  wire[46:0] twiddle4_1_16_imag;
  wire[46:0] T18861;
  wire[42:0] T18862;
  wire[42:0] T18863;
  wire[3:0] T18864;
  wire T18865;
  wire[46:0] T18866;
  wire[46:0] T18867;
  wire[46:0] twiddle4_1_17_imag;
  wire[46:0] T18868;
  wire[42:0] T18869;
  wire[42:0] T18870;
  wire[3:0] T18871;
  wire T18872;
  wire[46:0] T18873;
  wire[46:0] T18874;
  wire T18875;
  wire[46:0] T18876;
  wire[46:0] twiddle4_1_18_imag;
  wire[46:0] T18877;
  wire[42:0] T18878;
  wire[42:0] T18879;
  wire[3:0] T18880;
  wire T18881;
  wire[46:0] T18882;
  wire[46:0] T18883;
  wire[46:0] twiddle4_1_19_imag;
  wire[46:0] T18884;
  wire[42:0] T18885;
  wire[42:0] T18886;
  wire[3:0] T18887;
  wire T18888;
  wire[46:0] T18889;
  wire[46:0] T18890;
  wire T18891;
  wire T18892;
  wire[46:0] T18893;
  wire[46:0] T18894;
  wire[46:0] twiddle4_1_20_imag;
  wire[46:0] T18895;
  wire[42:0] T18896;
  wire[42:0] T18897;
  wire[3:0] T18898;
  wire T18899;
  wire[46:0] T18900;
  wire[46:0] T18901;
  wire[46:0] twiddle4_1_21_imag;
  wire[46:0] T18902;
  wire[43:0] T18903;
  wire[43:0] T18904;
  wire[2:0] T18905;
  wire T18906;
  wire[46:0] T18907;
  wire[46:0] T18908;
  wire T18909;
  wire[46:0] T18910;
  wire[46:0] twiddle4_1_22_imag;
  wire[46:0] T18911;
  wire[43:0] T18912;
  wire[43:0] T18913;
  wire[2:0] T18914;
  wire T18915;
  wire[46:0] T18916;
  wire[46:0] T18917;
  wire[46:0] twiddle4_1_23_imag;
  wire[46:0] T18918;
  wire[43:0] T18919;
  wire[43:0] T18920;
  wire[2:0] T18921;
  wire T18922;
  wire[46:0] T18923;
  wire[46:0] T18924;
  wire T18925;
  wire T18926;
  wire T18927;
  wire[46:0] T18928;
  wire[46:0] T18929;
  wire[46:0] T18930;
  wire[46:0] twiddle4_1_24_imag;
  wire[46:0] T18931;
  wire[43:0] T18932;
  wire[43:0] T18933;
  wire[2:0] T18934;
  wire T18935;
  wire[46:0] T18936;
  wire[46:0] T18937;
  wire[46:0] twiddle4_1_25_imag;
  wire[46:0] T18938;
  wire[43:0] T18939;
  wire[43:0] T18940;
  wire[2:0] T18941;
  wire T18942;
  wire[46:0] T18943;
  wire[46:0] T18944;
  wire T18945;
  wire[46:0] T18946;
  wire[46:0] twiddle4_1_26_imag;
  wire[46:0] T18947;
  wire[43:0] T18948;
  wire[43:0] T18949;
  wire[2:0] T18950;
  wire T18951;
  wire[46:0] T18952;
  wire[46:0] T18953;
  wire[46:0] twiddle4_1_27_imag;
  wire[46:0] T18954;
  wire[43:0] T18955;
  wire[43:0] T18956;
  wire[2:0] T18957;
  wire T18958;
  wire[46:0] T18959;
  wire[46:0] T18960;
  wire T18961;
  wire T18962;
  wire[46:0] T18963;
  wire[46:0] T18964;
  wire[46:0] twiddle4_1_28_imag;
  wire[46:0] T18965;
  wire[43:0] T18966;
  wire[43:0] T18967;
  wire[2:0] T18968;
  wire T18969;
  wire[46:0] T18970;
  wire[46:0] T18971;
  wire[46:0] twiddle4_1_29_imag;
  wire[46:0] T18972;
  wire[43:0] T18973;
  wire[43:0] T18974;
  wire[2:0] T18975;
  wire T18976;
  wire[46:0] T18977;
  wire[46:0] T18978;
  wire T18979;
  wire[46:0] T18980;
  wire[46:0] twiddle4_1_30_imag;
  wire[46:0] T18981;
  wire[43:0] T18982;
  wire[43:0] T18983;
  wire[2:0] T18984;
  wire T18985;
  wire[46:0] T18986;
  wire[46:0] T18987;
  wire[46:0] twiddle4_1_31_imag;
  wire[46:0] T18988;
  wire[43:0] T18989;
  wire[43:0] T18990;
  wire[2:0] T18991;
  wire T18992;
  wire[46:0] T18993;
  wire[46:0] T18994;
  wire T18995;
  wire T18996;
  wire T18997;
  wire T18998;
  wire T18999;
  wire T19000;
  wire[47:0] T19001;
  wire[46:0] T19002;
  wire[46:0] T19003;
  wire[46:0] T19004;
  wire[46:0] T19005;
  wire[46:0] T19006;
  wire[46:0] twiddle4_1_32_imag;
  wire[46:0] T19007;
  wire[43:0] T19008;
  wire[43:0] T19009;
  wire[2:0] T19010;
  wire T19011;
  wire[46:0] T19012;
  wire[46:0] T19013;
  wire[46:0] twiddle4_1_33_imag;
  wire[46:0] T19014;
  wire[43:0] T19015;
  wire[43:0] T19016;
  wire[2:0] T19017;
  wire T19018;
  wire[46:0] T19019;
  wire[46:0] T19020;
  wire T19021;
  wire[46:0] T19022;
  wire[46:0] twiddle4_1_34_imag;
  wire[46:0] T19023;
  wire[43:0] T19024;
  wire[43:0] T19025;
  wire[2:0] T19026;
  wire T19027;
  wire[46:0] T19028;
  wire[46:0] T19029;
  wire[46:0] twiddle4_1_35_imag;
  wire[46:0] T19030;
  wire[43:0] T19031;
  wire[43:0] T19032;
  wire[2:0] T19033;
  wire T19034;
  wire[46:0] T19035;
  wire[46:0] T19036;
  wire T19037;
  wire T19038;
  wire[46:0] T19039;
  wire[46:0] T19040;
  wire[46:0] twiddle4_1_36_imag;
  wire[46:0] T19041;
  wire[43:0] T19042;
  wire[43:0] T19043;
  wire[2:0] T19044;
  wire T19045;
  wire[46:0] T19046;
  wire[46:0] T19047;
  wire[46:0] twiddle4_1_37_imag;
  wire[46:0] T19048;
  wire[43:0] T19049;
  wire[43:0] T19050;
  wire[2:0] T19051;
  wire T19052;
  wire[46:0] T19053;
  wire[46:0] T19054;
  wire T19055;
  wire[46:0] T19056;
  wire[46:0] twiddle4_1_38_imag;
  wire[46:0] T19057;
  wire[43:0] T19058;
  wire[43:0] T19059;
  wire[2:0] T19060;
  wire T19061;
  wire[46:0] T19062;
  wire[46:0] T19063;
  wire[46:0] twiddle4_1_39_imag;
  wire[46:0] T19064;
  wire[43:0] T19065;
  wire[43:0] T19066;
  wire[2:0] T19067;
  wire T19068;
  wire[46:0] T19069;
  wire[46:0] T19070;
  wire T19071;
  wire T19072;
  wire T19073;
  wire[46:0] T19074;
  wire[46:0] T19075;
  wire[46:0] T19076;
  wire[46:0] twiddle4_1_40_imag;
  wire[46:0] T19077;
  wire[43:0] T19078;
  wire[43:0] T19079;
  wire[2:0] T19080;
  wire T19081;
  wire[46:0] T19082;
  wire[46:0] T19083;
  wire[46:0] twiddle4_1_41_imag;
  wire[46:0] T19084;
  wire[44:0] T19085;
  wire[44:0] T19086;
  wire[1:0] T19087;
  wire T19088;
  wire[46:0] T19089;
  wire[46:0] T19090;
  wire T19091;
  wire[46:0] T19092;
  wire[46:0] twiddle4_1_42_imag;
  wire[46:0] T19093;
  wire[44:0] T19094;
  wire[44:0] T19095;
  wire[1:0] T19096;
  wire T19097;
  wire[46:0] T19098;
  wire[46:0] T19099;
  wire[46:0] twiddle4_1_43_imag;
  wire[46:0] T19100;
  wire[44:0] T19101;
  wire[44:0] T19102;
  wire[1:0] T19103;
  wire T19104;
  wire[46:0] T19105;
  wire[46:0] T19106;
  wire T19107;
  wire T19108;
  wire[46:0] T19109;
  wire[46:0] T19110;
  wire[46:0] twiddle4_1_44_imag;
  wire[46:0] T19111;
  wire[44:0] T19112;
  wire[44:0] T19113;
  wire[1:0] T19114;
  wire T19115;
  wire[46:0] T19116;
  wire[46:0] T19117;
  wire[46:0] twiddle4_1_45_imag;
  wire[46:0] T19118;
  wire[44:0] T19119;
  wire[44:0] T19120;
  wire[1:0] T19121;
  wire T19122;
  wire[46:0] T19123;
  wire[46:0] T19124;
  wire T19125;
  wire[46:0] T19126;
  wire[46:0] twiddle4_1_46_imag;
  wire[46:0] T19127;
  wire[44:0] T19128;
  wire[44:0] T19129;
  wire[1:0] T19130;
  wire T19131;
  wire[46:0] T19132;
  wire[46:0] T19133;
  wire[46:0] twiddle4_1_47_imag;
  wire[46:0] T19134;
  wire[44:0] T19135;
  wire[44:0] T19136;
  wire[1:0] T19137;
  wire T19138;
  wire[46:0] T19139;
  wire[46:0] T19140;
  wire T19141;
  wire T19142;
  wire T19143;
  wire T19144;
  wire[46:0] T19145;
  wire[46:0] T19146;
  wire[46:0] T19147;
  wire[46:0] T19148;
  wire[46:0] twiddle4_1_48_imag;
  wire[46:0] T19149;
  wire[44:0] T19150;
  wire[44:0] T19151;
  wire[1:0] T19152;
  wire T19153;
  wire[46:0] T19154;
  wire[46:0] T19155;
  wire[46:0] twiddle4_1_49_imag;
  wire[46:0] T19156;
  wire[44:0] T19157;
  wire[44:0] T19158;
  wire[1:0] T19159;
  wire T19160;
  wire[46:0] T19161;
  wire[46:0] T19162;
  wire T19163;
  wire[46:0] T19164;
  wire[46:0] twiddle4_1_50_imag;
  wire[46:0] T19165;
  wire[44:0] T19166;
  wire[44:0] T19167;
  wire[1:0] T19168;
  wire T19169;
  wire[46:0] T19170;
  wire[46:0] T19171;
  wire[46:0] twiddle4_1_51_imag;
  wire[46:0] T19172;
  wire[44:0] T19173;
  wire[44:0] T19174;
  wire[1:0] T19175;
  wire T19176;
  wire[46:0] T19177;
  wire[46:0] T19178;
  wire T19179;
  wire T19180;
  wire[46:0] T19181;
  wire[46:0] T19182;
  wire[46:0] twiddle4_1_52_imag;
  wire[46:0] T19183;
  wire[44:0] T19184;
  wire[44:0] T19185;
  wire[1:0] T19186;
  wire T19187;
  wire[46:0] T19188;
  wire[46:0] T19189;
  wire[46:0] twiddle4_1_53_imag;
  wire[46:0] T19190;
  wire[44:0] T19191;
  wire[44:0] T19192;
  wire[1:0] T19193;
  wire T19194;
  wire[46:0] T19195;
  wire[46:0] T19196;
  wire T19197;
  wire[46:0] T19198;
  wire[46:0] twiddle4_1_54_imag;
  wire[46:0] T19199;
  wire[44:0] T19200;
  wire[44:0] T19201;
  wire[1:0] T19202;
  wire T19203;
  wire[46:0] T19204;
  wire[46:0] T19205;
  wire[46:0] twiddle4_1_55_imag;
  wire[46:0] T19206;
  wire[44:0] T19207;
  wire[44:0] T19208;
  wire[1:0] T19209;
  wire T19210;
  wire[46:0] T19211;
  wire[46:0] T19212;
  wire T19213;
  wire T19214;
  wire T19215;
  wire[46:0] T19216;
  wire[46:0] T19217;
  wire[46:0] T19218;
  wire[46:0] twiddle4_1_56_imag;
  wire[46:0] T19219;
  wire[44:0] T19220;
  wire[44:0] T19221;
  wire[1:0] T19222;
  wire T19223;
  wire[46:0] T19224;
  wire[46:0] T19225;
  wire[46:0] twiddle4_1_57_imag;
  wire[46:0] T19226;
  wire[44:0] T19227;
  wire[44:0] T19228;
  wire[1:0] T19229;
  wire T19230;
  wire[46:0] T19231;
  wire[46:0] T19232;
  wire T19233;
  wire[46:0] T19234;
  wire[46:0] twiddle4_1_58_imag;
  wire[46:0] T19235;
  wire[44:0] T19236;
  wire[44:0] T19237;
  wire[1:0] T19238;
  wire T19239;
  wire[46:0] T19240;
  wire[46:0] T19241;
  wire[46:0] twiddle4_1_59_imag;
  wire[46:0] T19242;
  wire[44:0] T19243;
  wire[44:0] T19244;
  wire[1:0] T19245;
  wire T19246;
  wire[46:0] T19247;
  wire[46:0] T19248;
  wire T19249;
  wire T19250;
  wire[46:0] T19251;
  wire[46:0] T19252;
  wire[46:0] twiddle4_1_60_imag;
  wire[46:0] T19253;
  wire[44:0] T19254;
  wire[44:0] T19255;
  wire[1:0] T19256;
  wire T19257;
  wire[46:0] T19258;
  wire[46:0] T19259;
  wire[46:0] twiddle4_1_61_imag;
  wire[46:0] T19260;
  wire[44:0] T19261;
  wire[44:0] T19262;
  wire[1:0] T19263;
  wire T19264;
  wire[46:0] T19265;
  wire[46:0] T19266;
  wire T19267;
  wire[46:0] T19268;
  wire[46:0] twiddle4_1_62_imag;
  wire[46:0] T19269;
  wire[44:0] T19270;
  wire[44:0] T19271;
  wire[1:0] T19272;
  wire T19273;
  wire[46:0] T19274;
  wire[46:0] T19275;
  wire[46:0] twiddle4_1_63_imag;
  wire[46:0] T19276;
  wire[44:0] T19277;
  wire[44:0] T19278;
  wire[1:0] T19279;
  wire T19280;
  wire[46:0] T19281;
  wire[46:0] T19282;
  wire T19283;
  wire T19284;
  wire T19285;
  wire T19286;
  wire T19287;
  wire T19288;
  wire T19289;
  wire[47:0] T19290;
  wire[46:0] T19291;
  wire[46:0] T19292;
  wire[46:0] T19293;
  wire[46:0] T19294;
  wire[46:0] T19295;
  wire[46:0] T19296;
  wire[46:0] twiddle4_1_64_imag;
  wire[46:0] T19297;
  wire[44:0] T19298;
  wire[44:0] T19299;
  wire[1:0] T19300;
  wire T19301;
  wire[46:0] T19302;
  wire[46:0] T19303;
  wire[46:0] twiddle4_1_65_imag;
  wire[46:0] T19304;
  wire[44:0] T19305;
  wire[44:0] T19306;
  wire[1:0] T19307;
  wire T19308;
  wire[46:0] T19309;
  wire[46:0] T19310;
  wire T19311;
  wire[46:0] T19312;
  wire[46:0] twiddle4_1_66_imag;
  wire[46:0] T19313;
  wire[44:0] T19314;
  wire[44:0] T19315;
  wire[1:0] T19316;
  wire T19317;
  wire[46:0] T19318;
  wire[46:0] T19319;
  wire[46:0] twiddle4_1_67_imag;
  wire[46:0] T19320;
  wire[44:0] T19321;
  wire[44:0] T19322;
  wire[1:0] T19323;
  wire T19324;
  wire[46:0] T19325;
  wire[46:0] T19326;
  wire T19327;
  wire T19328;
  wire[46:0] T19329;
  wire[46:0] T19330;
  wire[46:0] twiddle4_1_68_imag;
  wire[46:0] T19331;
  wire[44:0] T19332;
  wire[44:0] T19333;
  wire[1:0] T19334;
  wire T19335;
  wire[46:0] T19336;
  wire[46:0] T19337;
  wire[46:0] twiddle4_1_69_imag;
  wire[46:0] T19338;
  wire[44:0] T19339;
  wire[44:0] T19340;
  wire[1:0] T19341;
  wire T19342;
  wire[46:0] T19343;
  wire[46:0] T19344;
  wire T19345;
  wire[46:0] T19346;
  wire[46:0] twiddle4_1_70_imag;
  wire[46:0] T19347;
  wire[44:0] T19348;
  wire[44:0] T19349;
  wire[1:0] T19350;
  wire T19351;
  wire[46:0] T19352;
  wire[46:0] T19353;
  wire[46:0] twiddle4_1_71_imag;
  wire[46:0] T19354;
  wire[44:0] T19355;
  wire[44:0] T19356;
  wire[1:0] T19357;
  wire T19358;
  wire[46:0] T19359;
  wire[46:0] T19360;
  wire T19361;
  wire T19362;
  wire T19363;
  wire[46:0] T19364;
  wire[46:0] T19365;
  wire[46:0] T19366;
  wire[46:0] twiddle4_1_72_imag;
  wire[46:0] T19367;
  wire[44:0] T19368;
  wire[44:0] T19369;
  wire[1:0] T19370;
  wire T19371;
  wire[46:0] T19372;
  wire[46:0] T19373;
  wire[46:0] twiddle4_1_73_imag;
  wire[46:0] T19374;
  wire[44:0] T19375;
  wire[44:0] T19376;
  wire[1:0] T19377;
  wire T19378;
  wire[46:0] T19379;
  wire[46:0] T19380;
  wire T19381;
  wire[46:0] T19382;
  wire[46:0] twiddle4_1_74_imag;
  wire[46:0] T19383;
  wire[44:0] T19384;
  wire[44:0] T19385;
  wire[1:0] T19386;
  wire T19387;
  wire[46:0] T19388;
  wire[46:0] T19389;
  wire[46:0] twiddle4_1_75_imag;
  wire[46:0] T19390;
  wire[44:0] T19391;
  wire[44:0] T19392;
  wire[1:0] T19393;
  wire T19394;
  wire[46:0] T19395;
  wire[46:0] T19396;
  wire T19397;
  wire T19398;
  wire[46:0] T19399;
  wire[46:0] T19400;
  wire[46:0] twiddle4_1_76_imag;
  wire[46:0] T19401;
  wire[44:0] T19402;
  wire[44:0] T19403;
  wire[1:0] T19404;
  wire T19405;
  wire[46:0] T19406;
  wire[46:0] T19407;
  wire[46:0] twiddle4_1_77_imag;
  wire[46:0] T19408;
  wire[44:0] T19409;
  wire[44:0] T19410;
  wire[1:0] T19411;
  wire T19412;
  wire[46:0] T19413;
  wire[46:0] T19414;
  wire T19415;
  wire[46:0] T19416;
  wire[46:0] twiddle4_1_78_imag;
  wire[46:0] T19417;
  wire[44:0] T19418;
  wire[44:0] T19419;
  wire[1:0] T19420;
  wire T19421;
  wire[46:0] T19422;
  wire[46:0] T19423;
  wire[46:0] twiddle4_1_79_imag;
  wire[46:0] T19424;
  wire[44:0] T19425;
  wire[44:0] T19426;
  wire[1:0] T19427;
  wire T19428;
  wire[46:0] T19429;
  wire[46:0] T19430;
  wire T19431;
  wire T19432;
  wire T19433;
  wire T19434;
  wire[46:0] T19435;
  wire[46:0] T19436;
  wire[46:0] T19437;
  wire[46:0] T19438;
  wire[46:0] twiddle4_1_80_imag;
  wire[46:0] T19439;
  wire[44:0] T19440;
  wire[44:0] T19441;
  wire[1:0] T19442;
  wire T19443;
  wire[46:0] T19444;
  wire[46:0] T19445;
  wire[46:0] twiddle4_1_81_imag;
  wire[46:0] T19446;
  wire[44:0] T19447;
  wire[44:0] T19448;
  wire[1:0] T19449;
  wire T19450;
  wire[46:0] T19451;
  wire[46:0] T19452;
  wire T19453;
  wire[46:0] T19454;
  wire[46:0] twiddle4_1_82_imag;
  wire[46:0] T19455;
  wire[44:0] T19456;
  wire[44:0] T19457;
  wire[1:0] T19458;
  wire T19459;
  wire[46:0] T19460;
  wire[46:0] T19461;
  wire[46:0] twiddle4_1_83_imag;
  wire[46:0] T19462;
  wire[45:0] T19463;
  wire[45:0] T19464;
  wire T19465;
  wire[46:0] T19466;
  wire[46:0] T19467;
  wire T19468;
  wire T19469;
  wire[46:0] T19470;
  wire[46:0] T19471;
  wire[46:0] twiddle4_1_84_imag;
  wire[46:0] T19472;
  wire[45:0] T19473;
  wire[45:0] T19474;
  wire T19475;
  wire[46:0] T19476;
  wire[46:0] T19477;
  wire[46:0] twiddle4_1_85_imag;
  wire[46:0] T19478;
  wire[45:0] T19479;
  wire[45:0] T19480;
  wire T19481;
  wire[46:0] T19482;
  wire[46:0] T19483;
  wire T19484;
  wire[46:0] T19485;
  wire[46:0] twiddle4_1_86_imag;
  wire[46:0] T19486;
  wire[45:0] T19487;
  wire[45:0] T19488;
  wire T19489;
  wire[46:0] T19490;
  wire[46:0] T19491;
  wire[46:0] twiddle4_1_87_imag;
  wire[46:0] T19492;
  wire[45:0] T19493;
  wire[45:0] T19494;
  wire T19495;
  wire[46:0] T19496;
  wire[46:0] T19497;
  wire T19498;
  wire T19499;
  wire T19500;
  wire[46:0] T19501;
  wire[46:0] T19502;
  wire[46:0] T19503;
  wire[46:0] twiddle4_1_88_imag;
  wire[46:0] T19504;
  wire[45:0] T19505;
  wire[45:0] T19506;
  wire T19507;
  wire[46:0] T19508;
  wire[46:0] T19509;
  wire[46:0] twiddle4_1_89_imag;
  wire[46:0] T19510;
  wire[45:0] T19511;
  wire[45:0] T19512;
  wire T19513;
  wire[46:0] T19514;
  wire[46:0] T19515;
  wire T19516;
  wire[46:0] T19517;
  wire[46:0] twiddle4_1_90_imag;
  wire[46:0] T19518;
  wire[45:0] T19519;
  wire[45:0] T19520;
  wire T19521;
  wire[46:0] T19522;
  wire[46:0] T19523;
  wire[46:0] twiddle4_1_91_imag;
  wire[46:0] T19524;
  wire[45:0] T19525;
  wire[45:0] T19526;
  wire T19527;
  wire[46:0] T19528;
  wire[46:0] T19529;
  wire T19530;
  wire T19531;
  wire[46:0] T19532;
  wire[46:0] T19533;
  wire[46:0] twiddle4_1_92_imag;
  wire[46:0] T19534;
  wire[45:0] T19535;
  wire[45:0] T19536;
  wire T19537;
  wire[46:0] T19538;
  wire[46:0] T19539;
  wire[46:0] twiddle4_1_93_imag;
  wire[46:0] T19540;
  wire[45:0] T19541;
  wire[45:0] T19542;
  wire T19543;
  wire[46:0] T19544;
  wire[46:0] T19545;
  wire T19546;
  wire[46:0] T19547;
  wire[46:0] twiddle4_1_94_imag;
  wire[46:0] T19548;
  wire[45:0] T19549;
  wire[45:0] T19550;
  wire T19551;
  wire[46:0] T19552;
  wire[46:0] T19553;
  wire[46:0] twiddle4_1_95_imag;
  wire[46:0] T19554;
  wire[45:0] T19555;
  wire[45:0] T19556;
  wire T19557;
  wire[46:0] T19558;
  wire[46:0] T19559;
  wire T19560;
  wire T19561;
  wire T19562;
  wire T19563;
  wire T19564;
  wire[46:0] T19565;
  wire[46:0] T19566;
  wire[46:0] T19567;
  wire[46:0] T19568;
  wire[46:0] T19569;
  wire[46:0] twiddle4_1_96_imag;
  wire[46:0] T19570;
  wire[45:0] T19571;
  wire[45:0] T19572;
  wire T19573;
  wire[46:0] T19574;
  wire[46:0] T19575;
  wire[46:0] twiddle4_1_97_imag;
  wire[46:0] T19576;
  wire[45:0] T19577;
  wire[45:0] T19578;
  wire T19579;
  wire[46:0] T19580;
  wire[46:0] T19581;
  wire T19582;
  wire[46:0] T19583;
  wire[46:0] twiddle4_1_98_imag;
  wire[46:0] T19584;
  wire[45:0] T19585;
  wire[45:0] T19586;
  wire T19587;
  wire[46:0] T19588;
  wire[46:0] T19589;
  wire[46:0] twiddle4_1_99_imag;
  wire[46:0] T19590;
  wire[45:0] T19591;
  wire[45:0] T19592;
  wire T19593;
  wire[46:0] T19594;
  wire[46:0] T19595;
  wire T19596;
  wire T19597;
  wire[46:0] T19598;
  wire[46:0] T19599;
  wire[46:0] twiddle4_1_100_imag;
  wire[46:0] T19600;
  wire[45:0] T19601;
  wire[45:0] T19602;
  wire T19603;
  wire[46:0] T19604;
  wire[46:0] T19605;
  wire[46:0] twiddle4_1_101_imag;
  wire[46:0] T19606;
  wire[45:0] T19607;
  wire[45:0] T19608;
  wire T19609;
  wire[46:0] T19610;
  wire[46:0] T19611;
  wire T19612;
  wire[46:0] T19613;
  wire[46:0] twiddle4_1_102_imag;
  wire[46:0] T19614;
  wire[45:0] T19615;
  wire[45:0] T19616;
  wire T19617;
  wire[46:0] T19618;
  wire[46:0] T19619;
  wire[46:0] twiddle4_1_103_imag;
  wire[46:0] T19620;
  wire[45:0] T19621;
  wire[45:0] T19622;
  wire T19623;
  wire[46:0] T19624;
  wire[46:0] T19625;
  wire T19626;
  wire T19627;
  wire T19628;
  wire[46:0] T19629;
  wire[46:0] T19630;
  wire[46:0] T19631;
  wire[46:0] twiddle4_1_104_imag;
  wire[46:0] T19632;
  wire[45:0] T19633;
  wire[45:0] T19634;
  wire T19635;
  wire[46:0] T19636;
  wire[46:0] T19637;
  wire[46:0] twiddle4_1_105_imag;
  wire[46:0] T19638;
  wire[45:0] T19639;
  wire[45:0] T19640;
  wire T19641;
  wire[46:0] T19642;
  wire[46:0] T19643;
  wire T19644;
  wire[46:0] T19645;
  wire[46:0] twiddle4_1_106_imag;
  wire[46:0] T19646;
  wire[45:0] T19647;
  wire[45:0] T19648;
  wire T19649;
  wire[46:0] T19650;
  wire[46:0] T19651;
  wire[46:0] twiddle4_1_107_imag;
  wire[46:0] T19652;
  wire[45:0] T19653;
  wire[45:0] T19654;
  wire T19655;
  wire[46:0] T19656;
  wire[46:0] T19657;
  wire T19658;
  wire T19659;
  wire[46:0] T19660;
  wire[46:0] T19661;
  wire[46:0] twiddle4_1_108_imag;
  wire[46:0] T19662;
  wire[45:0] T19663;
  wire[45:0] T19664;
  wire T19665;
  wire[46:0] T19666;
  wire[46:0] T19667;
  wire[46:0] twiddle4_1_109_imag;
  wire[46:0] T19668;
  wire[45:0] T19669;
  wire[45:0] T19670;
  wire T19671;
  wire[46:0] T19672;
  wire[46:0] T19673;
  wire T19674;
  wire[46:0] T19675;
  wire[46:0] twiddle4_1_110_imag;
  wire[46:0] T19676;
  wire[45:0] T19677;
  wire[45:0] T19678;
  wire T19679;
  wire[46:0] T19680;
  wire[46:0] T19681;
  wire[46:0] twiddle4_1_111_imag;
  wire[46:0] T19682;
  wire[45:0] T19683;
  wire[45:0] T19684;
  wire T19685;
  wire[46:0] T19686;
  wire[46:0] T19687;
  wire T19688;
  wire T19689;
  wire T19690;
  wire T19691;
  wire[46:0] T19692;
  wire[46:0] T19693;
  wire[46:0] T19694;
  wire[46:0] T19695;
  wire[46:0] twiddle4_1_112_imag;
  wire[46:0] T19696;
  wire[45:0] T19697;
  wire[45:0] T19698;
  wire T19699;
  wire[46:0] T19700;
  wire[46:0] T19701;
  wire[46:0] twiddle4_1_113_imag;
  wire[46:0] T19702;
  wire[45:0] T19703;
  wire[45:0] T19704;
  wire T19705;
  wire[46:0] T19706;
  wire[46:0] T19707;
  wire T19708;
  wire[46:0] T19709;
  wire[46:0] twiddle4_1_114_imag;
  wire[46:0] T19710;
  wire[45:0] T19711;
  wire[45:0] T19712;
  wire T19713;
  wire[46:0] T19714;
  wire[46:0] T19715;
  wire[46:0] twiddle4_1_115_imag;
  wire[46:0] T19716;
  wire[45:0] T19717;
  wire[45:0] T19718;
  wire T19719;
  wire[46:0] T19720;
  wire[46:0] T19721;
  wire T19722;
  wire T19723;
  wire[46:0] T19724;
  wire[46:0] T19725;
  wire[46:0] twiddle4_1_116_imag;
  wire[46:0] T19726;
  wire[45:0] T19727;
  wire[45:0] T19728;
  wire T19729;
  wire[46:0] T19730;
  wire[46:0] T19731;
  wire[46:0] twiddle4_1_117_imag;
  wire[46:0] T19732;
  wire[45:0] T19733;
  wire[45:0] T19734;
  wire T19735;
  wire[46:0] T19736;
  wire[46:0] T19737;
  wire T19738;
  wire[46:0] T19739;
  wire[46:0] twiddle4_1_118_imag;
  wire[46:0] T19740;
  wire[45:0] T19741;
  wire[45:0] T19742;
  wire T19743;
  wire[46:0] T19744;
  wire[46:0] T19745;
  wire[46:0] twiddle4_1_119_imag;
  wire[46:0] T19746;
  wire[45:0] T19747;
  wire[45:0] T19748;
  wire T19749;
  wire[46:0] T19750;
  wire[46:0] T19751;
  wire T19752;
  wire T19753;
  wire T19754;
  wire[46:0] T19755;
  wire[46:0] T19756;
  wire[46:0] T19757;
  wire[46:0] twiddle4_1_120_imag;
  wire[46:0] T19758;
  wire[45:0] T19759;
  wire[45:0] T19760;
  wire T19761;
  wire[46:0] T19762;
  wire[46:0] T19763;
  wire[46:0] twiddle4_1_121_imag;
  wire[46:0] T19764;
  wire[45:0] T19765;
  wire[45:0] T19766;
  wire T19767;
  wire[46:0] T19768;
  wire[46:0] T19769;
  wire T19770;
  wire[46:0] T19771;
  wire[46:0] twiddle4_1_122_imag;
  wire[46:0] T19772;
  wire[45:0] T19773;
  wire[45:0] T19774;
  wire T19775;
  wire[46:0] T19776;
  wire[46:0] T19777;
  wire[46:0] twiddle4_1_123_imag;
  wire[46:0] T19778;
  wire[45:0] T19779;
  wire[45:0] T19780;
  wire T19781;
  wire[46:0] T19782;
  wire[46:0] T19783;
  wire T19784;
  wire T19785;
  wire[46:0] T19786;
  wire[46:0] T19787;
  wire[46:0] twiddle4_1_124_imag;
  wire[46:0] T19788;
  wire[45:0] T19789;
  wire[45:0] T19790;
  wire T19791;
  wire[46:0] T19792;
  wire[46:0] T19793;
  wire[46:0] twiddle4_1_125_imag;
  wire[46:0] T19794;
  wire[45:0] T19795;
  wire[45:0] T19796;
  wire T19797;
  wire[46:0] T19798;
  wire[46:0] T19799;
  wire T19800;
  wire[46:0] T19801;
  wire[46:0] twiddle4_1_126_imag;
  wire[46:0] T19802;
  wire[45:0] T19803;
  wire[45:0] T19804;
  wire T19805;
  wire[46:0] T19806;
  wire[46:0] T19807;
  wire[46:0] twiddle4_1_127_imag;
  wire[46:0] T19808;
  wire[45:0] T19809;
  wire[45:0] T19810;
  wire T19811;
  wire[46:0] T19812;
  wire[46:0] T19813;
  wire T19814;
  wire T19815;
  wire T19816;
  wire T19817;
  wire T19818;
  wire T19819;
  wire T19820;
  wire T19821;
  wire[47:0] T19822;
  wire[46:0] T19823;
  wire[46:0] T19824;
  wire[46:0] T19825;
  wire[46:0] T19826;
  wire[46:0] T19827;
  wire[46:0] T19828;
  wire[46:0] T19829;
  wire[46:0] twiddle4_1_128_imag;
  wire[46:0] T19830;
  wire[45:0] T19831;
  wire[45:0] T19832;
  wire T19833;
  wire[46:0] T19834;
  wire[46:0] T19835;
  wire[46:0] twiddle4_1_129_imag;
  wire[46:0] T19836;
  wire[45:0] T19837;
  wire[45:0] T19838;
  wire T19839;
  wire[46:0] T19840;
  wire[46:0] T19841;
  wire T19842;
  wire[46:0] T19843;
  wire[46:0] twiddle4_1_130_imag;
  wire[46:0] T19844;
  wire[45:0] T19845;
  wire[45:0] T19846;
  wire T19847;
  wire[46:0] T19848;
  wire[46:0] T19849;
  wire[46:0] twiddle4_1_131_imag;
  wire[46:0] T19850;
  wire[45:0] T19851;
  wire[45:0] T19852;
  wire T19853;
  wire[46:0] T19854;
  wire[46:0] T19855;
  wire T19856;
  wire T19857;
  wire[46:0] T19858;
  wire[46:0] T19859;
  wire[46:0] twiddle4_1_132_imag;
  wire[46:0] T19860;
  wire[45:0] T19861;
  wire[45:0] T19862;
  wire T19863;
  wire[46:0] T19864;
  wire[46:0] T19865;
  wire[46:0] twiddle4_1_133_imag;
  wire[46:0] T19866;
  wire[45:0] T19867;
  wire[45:0] T19868;
  wire T19869;
  wire[46:0] T19870;
  wire[46:0] T19871;
  wire T19872;
  wire[46:0] T19873;
  wire[46:0] twiddle4_1_134_imag;
  wire[46:0] T19874;
  wire[45:0] T19875;
  wire[45:0] T19876;
  wire T19877;
  wire[46:0] T19878;
  wire[46:0] T19879;
  wire[46:0] twiddle4_1_135_imag;
  wire[46:0] T19880;
  wire[45:0] T19881;
  wire[45:0] T19882;
  wire T19883;
  wire[46:0] T19884;
  wire[46:0] T19885;
  wire T19886;
  wire T19887;
  wire T19888;
  wire[46:0] T19889;
  wire[46:0] T19890;
  wire[46:0] T19891;
  wire[46:0] twiddle4_1_136_imag;
  wire[46:0] T19892;
  wire[45:0] T19893;
  wire[45:0] T19894;
  wire T19895;
  wire[46:0] T19896;
  wire[46:0] T19897;
  wire[46:0] twiddle4_1_137_imag;
  wire[46:0] T19898;
  wire[45:0] T19899;
  wire[45:0] T19900;
  wire T19901;
  wire[46:0] T19902;
  wire[46:0] T19903;
  wire T19904;
  wire[46:0] T19905;
  wire[46:0] twiddle4_1_138_imag;
  wire[46:0] T19906;
  wire[45:0] T19907;
  wire[45:0] T19908;
  wire T19909;
  wire[46:0] T19910;
  wire[46:0] T19911;
  wire[46:0] twiddle4_1_139_imag;
  wire[46:0] T19912;
  wire[45:0] T19913;
  wire[45:0] T19914;
  wire T19915;
  wire[46:0] T19916;
  wire[46:0] T19917;
  wire T19918;
  wire T19919;
  wire[46:0] T19920;
  wire[46:0] T19921;
  wire[46:0] twiddle4_1_140_imag;
  wire[46:0] T19922;
  wire[45:0] T19923;
  wire[45:0] T19924;
  wire T19925;
  wire[46:0] T19926;
  wire[46:0] T19927;
  wire[46:0] twiddle4_1_141_imag;
  wire[46:0] T19928;
  wire[45:0] T19929;
  wire[45:0] T19930;
  wire T19931;
  wire[46:0] T19932;
  wire[46:0] T19933;
  wire T19934;
  wire[46:0] T19935;
  wire[46:0] twiddle4_1_142_imag;
  wire[46:0] T19936;
  wire[45:0] T19937;
  wire[45:0] T19938;
  wire T19939;
  wire[46:0] T19940;
  wire[46:0] T19941;
  wire[46:0] twiddle4_1_143_imag;
  wire[46:0] T19942;
  wire[45:0] T19943;
  wire[45:0] T19944;
  wire T19945;
  wire[46:0] T19946;
  wire[46:0] T19947;
  wire T19948;
  wire T19949;
  wire T19950;
  wire T19951;
  wire[46:0] T19952;
  wire[46:0] T19953;
  wire[46:0] T19954;
  wire[46:0] T19955;
  wire[46:0] twiddle4_1_144_imag;
  wire[46:0] T19956;
  wire[45:0] T19957;
  wire[45:0] T19958;
  wire T19959;
  wire[46:0] T19960;
  wire[46:0] T19961;
  wire[46:0] twiddle4_1_145_imag;
  wire[46:0] T19962;
  wire[45:0] T19963;
  wire[45:0] T19964;
  wire T19965;
  wire[46:0] T19966;
  wire[46:0] T19967;
  wire T19968;
  wire[46:0] T19969;
  wire[46:0] twiddle4_1_146_imag;
  wire[46:0] T19970;
  wire[45:0] T19971;
  wire[45:0] T19972;
  wire T19973;
  wire[46:0] T19974;
  wire[46:0] T19975;
  wire[46:0] twiddle4_1_147_imag;
  wire[46:0] T19976;
  wire[45:0] T19977;
  wire[45:0] T19978;
  wire T19979;
  wire[46:0] T19980;
  wire[46:0] T19981;
  wire T19982;
  wire T19983;
  wire[46:0] T19984;
  wire[46:0] T19985;
  wire[46:0] twiddle4_1_148_imag;
  wire[46:0] T19986;
  wire[45:0] T19987;
  wire[45:0] T19988;
  wire T19989;
  wire[46:0] T19990;
  wire[46:0] T19991;
  wire[46:0] twiddle4_1_149_imag;
  wire[46:0] T19992;
  wire[45:0] T19993;
  wire[45:0] T19994;
  wire T19995;
  wire[46:0] T19996;
  wire[46:0] T19997;
  wire T19998;
  wire[46:0] T19999;
  wire[46:0] twiddle4_1_150_imag;
  wire[46:0] T20000;
  wire[45:0] T20001;
  wire[45:0] T20002;
  wire T20003;
  wire[46:0] T20004;
  wire[46:0] T20005;
  wire[46:0] twiddle4_1_151_imag;
  wire[46:0] T20006;
  wire[45:0] T20007;
  wire[45:0] T20008;
  wire T20009;
  wire[46:0] T20010;
  wire[46:0] T20011;
  wire T20012;
  wire T20013;
  wire T20014;
  wire[46:0] T20015;
  wire[46:0] T20016;
  wire[46:0] T20017;
  wire[46:0] twiddle4_1_152_imag;
  wire[46:0] T20018;
  wire[45:0] T20019;
  wire[45:0] T20020;
  wire T20021;
  wire[46:0] T20022;
  wire[46:0] T20023;
  wire[46:0] twiddle4_1_153_imag;
  wire[46:0] T20024;
  wire[45:0] T20025;
  wire[45:0] T20026;
  wire T20027;
  wire[46:0] T20028;
  wire[46:0] T20029;
  wire T20030;
  wire[46:0] T20031;
  wire[46:0] twiddle4_1_154_imag;
  wire[46:0] T20032;
  wire[45:0] T20033;
  wire[45:0] T20034;
  wire T20035;
  wire[46:0] T20036;
  wire[46:0] T20037;
  wire[46:0] twiddle4_1_155_imag;
  wire[46:0] T20038;
  wire[45:0] T20039;
  wire[45:0] T20040;
  wire T20041;
  wire[46:0] T20042;
  wire[46:0] T20043;
  wire T20044;
  wire T20045;
  wire[46:0] T20046;
  wire[46:0] T20047;
  wire[46:0] twiddle4_1_156_imag;
  wire[46:0] T20048;
  wire[45:0] T20049;
  wire[45:0] T20050;
  wire T20051;
  wire[46:0] T20052;
  wire[46:0] T20053;
  wire[46:0] twiddle4_1_157_imag;
  wire[46:0] T20054;
  wire[45:0] T20055;
  wire[45:0] T20056;
  wire T20057;
  wire[46:0] T20058;
  wire[46:0] T20059;
  wire T20060;
  wire[46:0] T20061;
  wire[46:0] twiddle4_1_158_imag;
  wire[46:0] T20062;
  wire[45:0] T20063;
  wire[45:0] T20064;
  wire T20065;
  wire[46:0] T20066;
  wire[46:0] T20067;
  wire[46:0] twiddle4_1_159_imag;
  wire[46:0] T20068;
  wire[45:0] T20069;
  wire[45:0] T20070;
  wire T20071;
  wire[46:0] T20072;
  wire[46:0] T20073;
  wire T20074;
  wire T20075;
  wire T20076;
  wire T20077;
  wire T20078;
  wire[46:0] T20079;
  wire[46:0] T20080;
  wire[46:0] T20081;
  wire[46:0] T20082;
  wire[46:0] T20083;
  wire[46:0] twiddle4_1_160_imag;
  wire[46:0] T20084;
  wire[45:0] T20085;
  wire[45:0] T20086;
  wire T20087;
  wire[46:0] T20088;
  wire[46:0] T20089;
  wire[46:0] twiddle4_1_161_imag;
  wire[46:0] T20090;
  wire[45:0] T20091;
  wire[45:0] T20092;
  wire T20093;
  wire[46:0] T20094;
  wire[46:0] T20095;
  wire T20096;
  wire[46:0] T20097;
  wire[46:0] twiddle4_1_162_imag;
  wire[46:0] T20098;
  wire[45:0] T20099;
  wire[45:0] T20100;
  wire T20101;
  wire[46:0] T20102;
  wire[46:0] T20103;
  wire[46:0] twiddle4_1_163_imag;
  wire[46:0] T20104;
  wire[45:0] T20105;
  wire[45:0] T20106;
  wire T20107;
  wire[46:0] T20108;
  wire[46:0] T20109;
  wire T20110;
  wire T20111;
  wire[46:0] T20112;
  wire[46:0] T20113;
  wire[46:0] twiddle4_1_164_imag;
  wire[46:0] T20114;
  wire[45:0] T20115;
  wire[45:0] T20116;
  wire T20117;
  wire[46:0] T20118;
  wire[46:0] T20119;
  wire[46:0] twiddle4_1_165_imag;
  wire[46:0] T20120;
  wire[45:0] T20121;
  wire[45:0] T20122;
  wire T20123;
  wire[46:0] T20124;
  wire[46:0] T20125;
  wire T20126;
  wire[46:0] T20127;
  wire[46:0] twiddle4_1_166_imag;
  wire[46:0] T20128;
  wire[45:0] T20129;
  wire[45:0] T20130;
  wire T20131;
  wire[46:0] T20132;
  wire[46:0] T20133;
  wire[46:0] twiddle4_1_167_imag;
  wire[46:0] T20134;
  wire[45:0] T20135;
  wire[45:0] T20136;
  wire T20137;
  wire[46:0] T20138;
  wire[46:0] T20139;
  wire T20140;
  wire T20141;
  wire T20142;
  wire[46:0] T20143;
  wire[46:0] T20144;
  wire[46:0] T20145;
  wire[46:0] twiddle4_1_168_imag;
  wire[46:0] T20146;
  wire[45:0] T20147;
  wire[45:0] T20148;
  wire T20149;
  wire[46:0] T20150;
  wire[46:0] T20151;
  wire[46:0] twiddle4_1_169_imag;
  wire[46:0] T20152;
  wire[45:0] T20153;
  wire[45:0] T20154;
  wire T20155;
  wire[46:0] T20156;
  wire[46:0] T20157;
  wire T20158;
  wire[46:0] T20159;
  wire[46:0] twiddle4_1_170_imag;
  wire[46:0] T20160;
  wire[45:0] T20161;
  wire[45:0] T20162;
  wire T20163;
  wire[46:0] T20164;
  wire[46:0] T20165;
  wire[46:0] twiddle4_1_171_imag;
  wire[46:0] T20166;
  wire[46:0] T20167;
  wire[46:0] T20168;
  wire[46:0] T20169;
  wire T20170;
  wire T20171;
  wire[46:0] T20172;
  wire[46:0] T20173;
  wire[46:0] twiddle4_1_172_imag;
  wire[46:0] T20174;
  wire[46:0] T20175;
  wire[46:0] T20176;
  wire[46:0] T20177;
  wire[46:0] twiddle4_1_173_imag;
  wire[46:0] T20178;
  wire[46:0] T20179;
  wire[46:0] T20180;
  wire[46:0] T20181;
  wire T20182;
  wire[46:0] T20183;
  wire[46:0] twiddle4_1_174_imag;
  wire[46:0] T20184;
  wire[46:0] T20185;
  wire[46:0] T20186;
  wire[46:0] T20187;
  wire[46:0] twiddle4_1_175_imag;
  wire[46:0] T20188;
  wire[46:0] T20189;
  wire[46:0] T20190;
  wire[46:0] T20191;
  wire T20192;
  wire T20193;
  wire T20194;
  wire T20195;
  wire[46:0] T20196;
  wire[46:0] T20197;
  wire[46:0] T20198;
  wire[46:0] T20199;
  wire[46:0] twiddle4_1_176_imag;
  wire[46:0] T20200;
  wire[46:0] T20201;
  wire[46:0] T20202;
  wire[46:0] T20203;
  wire[46:0] twiddle4_1_177_imag;
  wire[46:0] T20204;
  wire[46:0] T20205;
  wire[46:0] T20206;
  wire[46:0] T20207;
  wire T20208;
  wire[46:0] T20209;
  wire[46:0] twiddle4_1_178_imag;
  wire[46:0] T20210;
  wire[46:0] T20211;
  wire[46:0] T20212;
  wire[46:0] T20213;
  wire[46:0] twiddle4_1_179_imag;
  wire[46:0] T20214;
  wire[46:0] T20215;
  wire[46:0] T20216;
  wire[46:0] T20217;
  wire T20218;
  wire T20219;
  wire[46:0] T20220;
  wire[46:0] T20221;
  wire[46:0] twiddle4_1_180_imag;
  wire[46:0] T20222;
  wire[46:0] T20223;
  wire[46:0] T20224;
  wire[46:0] T20225;
  wire[46:0] twiddle4_1_181_imag;
  wire[46:0] T20226;
  wire[46:0] T20227;
  wire[46:0] T20228;
  wire[46:0] T20229;
  wire T20230;
  wire[46:0] T20231;
  wire[46:0] twiddle4_1_182_imag;
  wire[46:0] T20232;
  wire[46:0] T20233;
  wire[46:0] T20234;
  wire[46:0] T20235;
  wire[46:0] twiddle4_1_183_imag;
  wire[46:0] T20236;
  wire[46:0] T20237;
  wire[46:0] T20238;
  wire[46:0] T20239;
  wire T20240;
  wire T20241;
  wire T20242;
  wire[46:0] T20243;
  wire[46:0] T20244;
  wire[46:0] T20245;
  wire[46:0] twiddle4_1_184_imag;
  wire[46:0] T20246;
  wire[46:0] T20247;
  wire[46:0] T20248;
  wire[46:0] T20249;
  wire[46:0] twiddle4_1_185_imag;
  wire[46:0] T20250;
  wire[46:0] T20251;
  wire[46:0] T20252;
  wire[46:0] T20253;
  wire T20254;
  wire[46:0] T20255;
  wire[46:0] twiddle4_1_186_imag;
  wire[46:0] T20256;
  wire[46:0] T20257;
  wire[46:0] T20258;
  wire[46:0] T20259;
  wire[46:0] twiddle4_1_187_imag;
  wire[46:0] T20260;
  wire[46:0] T20261;
  wire[46:0] T20262;
  wire[46:0] T20263;
  wire T20264;
  wire T20265;
  wire[46:0] T20266;
  wire[46:0] T20267;
  wire[46:0] twiddle4_1_188_imag;
  wire[46:0] T20268;
  wire[46:0] T20269;
  wire[46:0] T20270;
  wire[46:0] T20271;
  wire[46:0] twiddle4_1_189_imag;
  wire[46:0] T20272;
  wire[46:0] T20273;
  wire[46:0] T20274;
  wire[46:0] T20275;
  wire T20276;
  wire[46:0] T20277;
  wire[46:0] twiddle4_1_190_imag;
  wire[46:0] T20278;
  wire[46:0] T20279;
  wire[46:0] T20280;
  wire[46:0] T20281;
  wire[46:0] twiddle4_1_191_imag;
  wire[46:0] T20282;
  wire[46:0] T20283;
  wire[46:0] T20284;
  wire[46:0] T20285;
  wire T20286;
  wire T20287;
  wire T20288;
  wire T20289;
  wire T20290;
  wire T20291;
  wire[46:0] T20292;
  wire[46:0] T20293;
  wire[46:0] T20294;
  wire[46:0] T20295;
  wire[46:0] T20296;
  wire[46:0] T20297;
  wire[46:0] twiddle4_1_192_imag;
  wire[46:0] T20298;
  wire[46:0] T20299;
  wire[46:0] T20300;
  wire[46:0] T20301;
  wire[46:0] twiddle4_1_193_imag;
  wire[46:0] T20302;
  wire[46:0] T20303;
  wire[46:0] T20304;
  wire[46:0] T20305;
  wire T20306;
  wire[46:0] T20307;
  wire[46:0] twiddle4_1_194_imag;
  wire[46:0] T20308;
  wire[46:0] T20309;
  wire[46:0] T20310;
  wire[46:0] T20311;
  wire[46:0] twiddle4_1_195_imag;
  wire[46:0] T20312;
  wire[46:0] T20313;
  wire[46:0] T20314;
  wire[46:0] T20315;
  wire T20316;
  wire T20317;
  wire[46:0] T20318;
  wire[46:0] T20319;
  wire[46:0] twiddle4_1_196_imag;
  wire[46:0] T20320;
  wire[46:0] T20321;
  wire[46:0] T20322;
  wire[46:0] T20323;
  wire[46:0] twiddle4_1_197_imag;
  wire[46:0] T20324;
  wire[46:0] T20325;
  wire[46:0] T20326;
  wire[46:0] T20327;
  wire T20328;
  wire[46:0] T20329;
  wire[46:0] twiddle4_1_198_imag;
  wire[46:0] T20330;
  wire[46:0] T20331;
  wire[46:0] T20332;
  wire[46:0] T20333;
  wire[46:0] twiddle4_1_199_imag;
  wire[46:0] T20334;
  wire[46:0] T20335;
  wire[46:0] T20336;
  wire[46:0] T20337;
  wire T20338;
  wire T20339;
  wire T20340;
  wire[46:0] T20341;
  wire[46:0] T20342;
  wire[46:0] T20343;
  wire[46:0] twiddle4_1_200_imag;
  wire[46:0] T20344;
  wire[46:0] T20345;
  wire[46:0] T20346;
  wire[46:0] T20347;
  wire[46:0] twiddle4_1_201_imag;
  wire[46:0] T20348;
  wire[46:0] T20349;
  wire[46:0] T20350;
  wire[46:0] T20351;
  wire T20352;
  wire[46:0] T20353;
  wire[46:0] twiddle4_1_202_imag;
  wire[46:0] T20354;
  wire[46:0] T20355;
  wire[46:0] T20356;
  wire[46:0] T20357;
  wire[46:0] twiddle4_1_203_imag;
  wire[46:0] T20358;
  wire[46:0] T20359;
  wire[46:0] T20360;
  wire[46:0] T20361;
  wire T20362;
  wire T20363;
  wire[46:0] T20364;
  wire[46:0] T20365;
  wire[46:0] twiddle4_1_204_imag;
  wire[46:0] T20366;
  wire[46:0] T20367;
  wire[46:0] T20368;
  wire[46:0] T20369;
  wire[46:0] twiddle4_1_205_imag;
  wire[46:0] T20370;
  wire[46:0] T20371;
  wire[46:0] T20372;
  wire[46:0] T20373;
  wire T20374;
  wire[46:0] T20375;
  wire[46:0] twiddle4_1_206_imag;
  wire[46:0] T20376;
  wire[46:0] T20377;
  wire[46:0] T20378;
  wire[46:0] T20379;
  wire[46:0] twiddle4_1_207_imag;
  wire[46:0] T20380;
  wire[46:0] T20381;
  wire[46:0] T20382;
  wire[46:0] T20383;
  wire T20384;
  wire T20385;
  wire T20386;
  wire T20387;
  wire[46:0] T20388;
  wire[46:0] T20389;
  wire[46:0] T20390;
  wire[46:0] T20391;
  wire[46:0] twiddle4_1_208_imag;
  wire[46:0] T20392;
  wire[46:0] T20393;
  wire[46:0] T20394;
  wire[46:0] T20395;
  wire[46:0] twiddle4_1_209_imag;
  wire[46:0] T20396;
  wire[46:0] T20397;
  wire[46:0] T20398;
  wire[46:0] T20399;
  wire T20400;
  wire[46:0] T20401;
  wire[46:0] twiddle4_1_210_imag;
  wire[46:0] T20402;
  wire[46:0] T20403;
  wire[46:0] T20404;
  wire[46:0] T20405;
  wire[46:0] twiddle4_1_211_imag;
  wire[46:0] T20406;
  wire[46:0] T20407;
  wire[46:0] T20408;
  wire[46:0] T20409;
  wire T20410;
  wire T20411;
  wire[46:0] T20412;
  wire[46:0] T20413;
  wire[46:0] twiddle4_1_212_imag;
  wire[46:0] T20414;
  wire[46:0] T20415;
  wire[46:0] T20416;
  wire[46:0] T20417;
  wire[46:0] twiddle4_1_213_imag;
  wire[46:0] T20418;
  wire[46:0] T20419;
  wire[46:0] T20420;
  wire[46:0] T20421;
  wire T20422;
  wire[46:0] T20423;
  wire[46:0] twiddle4_1_214_imag;
  wire[46:0] T20424;
  wire[46:0] T20425;
  wire[46:0] T20426;
  wire[46:0] T20427;
  wire[46:0] twiddle4_1_215_imag;
  wire[46:0] T20428;
  wire[46:0] T20429;
  wire[46:0] T20430;
  wire[46:0] T20431;
  wire T20432;
  wire T20433;
  wire T20434;
  wire[46:0] T20435;
  wire[46:0] T20436;
  wire[46:0] T20437;
  wire[46:0] twiddle4_1_216_imag;
  wire[46:0] T20438;
  wire[46:0] T20439;
  wire[46:0] T20440;
  wire[46:0] T20441;
  wire[46:0] twiddle4_1_217_imag;
  wire[46:0] T20442;
  wire[46:0] T20443;
  wire[46:0] T20444;
  wire[46:0] T20445;
  wire T20446;
  wire[46:0] T20447;
  wire[46:0] twiddle4_1_218_imag;
  wire[46:0] T20448;
  wire[46:0] T20449;
  wire[46:0] T20450;
  wire[46:0] T20451;
  wire[46:0] twiddle4_1_219_imag;
  wire[46:0] T20452;
  wire[46:0] T20453;
  wire[46:0] T20454;
  wire[46:0] T20455;
  wire T20456;
  wire T20457;
  wire[46:0] T20458;
  wire[46:0] T20459;
  wire[46:0] twiddle4_1_220_imag;
  wire[46:0] T20460;
  wire[46:0] T20461;
  wire[46:0] T20462;
  wire[46:0] T20463;
  wire[46:0] twiddle4_1_221_imag;
  wire[46:0] T20464;
  wire[46:0] T20465;
  wire[46:0] T20466;
  wire[46:0] T20467;
  wire T20468;
  wire[46:0] T20469;
  wire[46:0] twiddle4_1_222_imag;
  wire[46:0] T20470;
  wire[46:0] T20471;
  wire[46:0] T20472;
  wire[46:0] T20473;
  wire[46:0] twiddle4_1_223_imag;
  wire[46:0] T20474;
  wire[46:0] T20475;
  wire[46:0] T20476;
  wire[46:0] T20477;
  wire T20478;
  wire T20479;
  wire T20480;
  wire T20481;
  wire T20482;
  wire[46:0] T20483;
  wire[46:0] T20484;
  wire[46:0] T20485;
  wire[46:0] T20486;
  wire[46:0] T20487;
  wire[46:0] twiddle4_1_224_imag;
  wire[46:0] T20488;
  wire[46:0] T20489;
  wire[46:0] T20490;
  wire[46:0] T20491;
  wire[46:0] twiddle4_1_225_imag;
  wire[46:0] T20492;
  wire[46:0] T20493;
  wire[46:0] T20494;
  wire[46:0] T20495;
  wire T20496;
  wire[46:0] T20497;
  wire[46:0] twiddle4_1_226_imag;
  wire[46:0] T20498;
  wire[46:0] T20499;
  wire[46:0] T20500;
  wire[46:0] T20501;
  wire[46:0] twiddle4_1_227_imag;
  wire[46:0] T20502;
  wire[46:0] T20503;
  wire[46:0] T20504;
  wire[46:0] T20505;
  wire T20506;
  wire T20507;
  wire[46:0] T20508;
  wire[46:0] T20509;
  wire[46:0] twiddle4_1_228_imag;
  wire[46:0] T20510;
  wire[46:0] T20511;
  wire[46:0] T20512;
  wire[46:0] T20513;
  wire[46:0] twiddle4_1_229_imag;
  wire[46:0] T20514;
  wire[46:0] T20515;
  wire[46:0] T20516;
  wire[46:0] T20517;
  wire T20518;
  wire[46:0] T20519;
  wire[46:0] twiddle4_1_230_imag;
  wire[46:0] T20520;
  wire[46:0] T20521;
  wire[46:0] T20522;
  wire[46:0] T20523;
  wire[46:0] twiddle4_1_231_imag;
  wire[46:0] T20524;
  wire[46:0] T20525;
  wire[46:0] T20526;
  wire[46:0] T20527;
  wire T20528;
  wire T20529;
  wire T20530;
  wire[46:0] T20531;
  wire[46:0] T20532;
  wire[46:0] T20533;
  wire[46:0] twiddle4_1_232_imag;
  wire[46:0] T20534;
  wire[46:0] T20535;
  wire[46:0] T20536;
  wire[46:0] T20537;
  wire[46:0] twiddle4_1_233_imag;
  wire[46:0] T20538;
  wire[46:0] T20539;
  wire[46:0] T20540;
  wire[46:0] T20541;
  wire T20542;
  wire[46:0] T20543;
  wire[46:0] twiddle4_1_234_imag;
  wire[46:0] T20544;
  wire[46:0] T20545;
  wire[46:0] T20546;
  wire[46:0] T20547;
  wire[46:0] twiddle4_1_235_imag;
  wire[46:0] T20548;
  wire[46:0] T20549;
  wire[46:0] T20550;
  wire[46:0] T20551;
  wire T20552;
  wire T20553;
  wire[46:0] T20554;
  wire[46:0] T20555;
  wire[46:0] twiddle4_1_236_imag;
  wire[46:0] T20556;
  wire[46:0] T20557;
  wire[46:0] T20558;
  wire[46:0] T20559;
  wire[46:0] twiddle4_1_237_imag;
  wire[46:0] T20560;
  wire[46:0] T20561;
  wire[46:0] T20562;
  wire[46:0] T20563;
  wire T20564;
  wire[46:0] T20565;
  wire[46:0] twiddle4_1_238_imag;
  wire[46:0] T20566;
  wire[46:0] T20567;
  wire[46:0] T20568;
  wire[46:0] T20569;
  wire[46:0] twiddle4_1_239_imag;
  wire[46:0] T20570;
  wire[46:0] T20571;
  wire[46:0] T20572;
  wire[46:0] T20573;
  wire T20574;
  wire T20575;
  wire T20576;
  wire T20577;
  wire[46:0] T20578;
  wire[46:0] T20579;
  wire[46:0] T20580;
  wire[46:0] T20581;
  wire[46:0] twiddle4_1_240_imag;
  wire[46:0] T20582;
  wire[46:0] T20583;
  wire[46:0] T20584;
  wire[46:0] T20585;
  wire[46:0] twiddle4_1_241_imag;
  wire[46:0] T20586;
  wire[46:0] T20587;
  wire[46:0] T20588;
  wire[46:0] T20589;
  wire T20590;
  wire[46:0] T20591;
  wire[46:0] twiddle4_1_242_imag;
  wire[46:0] T20592;
  wire[46:0] T20593;
  wire[46:0] T20594;
  wire[46:0] T20595;
  wire[46:0] twiddle4_1_243_imag;
  wire[46:0] T20596;
  wire[46:0] T20597;
  wire[46:0] T20598;
  wire[46:0] T20599;
  wire T20600;
  wire T20601;
  wire[46:0] T20602;
  wire[46:0] T20603;
  wire[46:0] twiddle4_1_244_imag;
  wire[46:0] T20604;
  wire[46:0] T20605;
  wire[46:0] T20606;
  wire[46:0] T20607;
  wire[46:0] twiddle4_1_245_imag;
  wire[46:0] T20608;
  wire[46:0] T20609;
  wire[46:0] T20610;
  wire[46:0] T20611;
  wire T20612;
  wire[46:0] T20613;
  wire[46:0] twiddle4_1_246_imag;
  wire[46:0] T20614;
  wire[46:0] T20615;
  wire[46:0] T20616;
  wire[46:0] T20617;
  wire[46:0] twiddle4_1_247_imag;
  wire[46:0] T20618;
  wire[46:0] T20619;
  wire[46:0] T20620;
  wire[46:0] T20621;
  wire T20622;
  wire T20623;
  wire T20624;
  wire[46:0] T20625;
  wire[46:0] T20626;
  wire[46:0] T20627;
  wire[46:0] twiddle4_1_248_imag;
  wire[46:0] T20628;
  wire[46:0] T20629;
  wire[46:0] T20630;
  wire[46:0] T20631;
  wire[46:0] twiddle4_1_249_imag;
  wire[46:0] T20632;
  wire[46:0] T20633;
  wire[46:0] T20634;
  wire[46:0] T20635;
  wire T20636;
  wire[46:0] T20637;
  wire[46:0] twiddle4_1_250_imag;
  wire[46:0] T20638;
  wire[46:0] T20639;
  wire[46:0] T20640;
  wire[46:0] T20641;
  wire[46:0] twiddle4_1_251_imag;
  wire[46:0] T20642;
  wire[46:0] T20643;
  wire[46:0] T20644;
  wire[46:0] T20645;
  wire T20646;
  wire T20647;
  wire[46:0] T20648;
  wire[46:0] T20649;
  wire[46:0] twiddle4_1_252_imag;
  wire[46:0] T20650;
  wire[46:0] T20651;
  wire[46:0] T20652;
  wire[46:0] T20653;
  wire[46:0] twiddle4_1_253_imag;
  wire[46:0] T20654;
  wire[46:0] T20655;
  wire[46:0] T20656;
  wire[46:0] T20657;
  wire T20658;
  wire[46:0] T20659;
  wire[46:0] twiddle4_1_254_imag;
  wire[46:0] T20660;
  wire[46:0] T20661;
  wire[46:0] T20662;
  wire[46:0] T20663;
  wire[46:0] twiddle4_1_255_imag;
  wire[46:0] T20664;
  wire[46:0] T20665;
  wire[46:0] T20666;
  wire[46:0] T20667;
  wire T20668;
  wire T20669;
  wire T20670;
  wire T20671;
  wire T20672;
  wire T20673;
  wire T20674;
  wire T20675;
  wire T20676;
  wire[47:0] T20677;
  wire[46:0] T20678;
  wire[46:0] T20679;
  wire[46:0] T20680;
  wire[46:0] T20681;
  wire[46:0] T20682;
  wire[46:0] T20683;
  wire[46:0] T20684;
  wire[46:0] T20685;
  wire[46:0] twiddle4_1_256_imag;
  wire[46:0] T20686;
  wire[46:0] T20687;
  wire[46:0] T20688;
  wire[46:0] T20689;
  wire[46:0] twiddle4_1_257_imag;
  wire[46:0] T20690;
  wire[46:0] T20691;
  wire[46:0] T20692;
  wire[46:0] T20693;
  wire T20694;
  wire[46:0] T20695;
  wire[46:0] twiddle4_1_258_imag;
  wire[46:0] T20696;
  wire[46:0] T20697;
  wire[46:0] T20698;
  wire[46:0] T20699;
  wire[46:0] twiddle4_1_259_imag;
  wire[46:0] T20700;
  wire[46:0] T20701;
  wire[46:0] T20702;
  wire[46:0] T20703;
  wire T20704;
  wire T20705;
  wire[46:0] T20706;
  wire[46:0] T20707;
  wire[46:0] twiddle4_1_260_imag;
  wire[46:0] T20708;
  wire[46:0] T20709;
  wire[46:0] T20710;
  wire[46:0] T20711;
  wire[46:0] twiddle4_1_261_imag;
  wire[46:0] T20712;
  wire[46:0] T20713;
  wire[46:0] T20714;
  wire[46:0] T20715;
  wire T20716;
  wire[46:0] T20717;
  wire[46:0] twiddle4_1_262_imag;
  wire[46:0] T20718;
  wire[46:0] T20719;
  wire[46:0] T20720;
  wire[46:0] T20721;
  wire[46:0] twiddle4_1_263_imag;
  wire[46:0] T20722;
  wire[46:0] T20723;
  wire[46:0] T20724;
  wire[46:0] T20725;
  wire T20726;
  wire T20727;
  wire T20728;
  wire[46:0] T20729;
  wire[46:0] T20730;
  wire[46:0] T20731;
  wire[46:0] twiddle4_1_264_imag;
  wire[46:0] T20732;
  wire[46:0] T20733;
  wire[46:0] T20734;
  wire[46:0] T20735;
  wire[46:0] twiddle4_1_265_imag;
  wire[46:0] T20736;
  wire[46:0] T20737;
  wire[46:0] T20738;
  wire[46:0] T20739;
  wire T20740;
  wire[46:0] T20741;
  wire[46:0] twiddle4_1_266_imag;
  wire[46:0] T20742;
  wire[46:0] T20743;
  wire[46:0] T20744;
  wire[46:0] T20745;
  wire[46:0] twiddle4_1_267_imag;
  wire[46:0] T20746;
  wire[46:0] T20747;
  wire[46:0] T20748;
  wire[46:0] T20749;
  wire T20750;
  wire T20751;
  wire[46:0] T20752;
  wire[46:0] T20753;
  wire[46:0] twiddle4_1_268_imag;
  wire[46:0] T20754;
  wire[46:0] T20755;
  wire[46:0] T20756;
  wire[46:0] T20757;
  wire[46:0] twiddle4_1_269_imag;
  wire[46:0] T20758;
  wire[46:0] T20759;
  wire[46:0] T20760;
  wire[46:0] T20761;
  wire T20762;
  wire[46:0] T20763;
  wire[46:0] twiddle4_1_270_imag;
  wire[46:0] T20764;
  wire[46:0] T20765;
  wire[46:0] T20766;
  wire[46:0] T20767;
  wire[46:0] twiddle4_1_271_imag;
  wire[46:0] T20768;
  wire[46:0] T20769;
  wire[46:0] T20770;
  wire[46:0] T20771;
  wire T20772;
  wire T20773;
  wire T20774;
  wire T20775;
  wire[46:0] T20776;
  wire[46:0] T20777;
  wire[46:0] T20778;
  wire[46:0] T20779;
  wire[46:0] twiddle4_1_272_imag;
  wire[46:0] T20780;
  wire[46:0] T20781;
  wire[46:0] T20782;
  wire[46:0] T20783;
  wire[46:0] twiddle4_1_273_imag;
  wire[46:0] T20784;
  wire[46:0] T20785;
  wire[46:0] T20786;
  wire[46:0] T20787;
  wire T20788;
  wire[46:0] T20789;
  wire[46:0] twiddle4_1_274_imag;
  wire[46:0] T20790;
  wire[46:0] T20791;
  wire[46:0] T20792;
  wire[46:0] T20793;
  wire[46:0] twiddle4_1_275_imag;
  wire[46:0] T20794;
  wire[46:0] T20795;
  wire[46:0] T20796;
  wire[46:0] T20797;
  wire T20798;
  wire T20799;
  wire[46:0] T20800;
  wire[46:0] T20801;
  wire[46:0] twiddle4_1_276_imag;
  wire[46:0] T20802;
  wire[46:0] T20803;
  wire[46:0] T20804;
  wire[46:0] T20805;
  wire[46:0] twiddle4_1_277_imag;
  wire[46:0] T20806;
  wire[46:0] T20807;
  wire[46:0] T20808;
  wire[46:0] T20809;
  wire T20810;
  wire[46:0] T20811;
  wire[46:0] twiddle4_1_278_imag;
  wire[46:0] T20812;
  wire[46:0] T20813;
  wire[46:0] T20814;
  wire[46:0] T20815;
  wire[46:0] twiddle4_1_279_imag;
  wire[46:0] T20816;
  wire[46:0] T20817;
  wire[46:0] T20818;
  wire[46:0] T20819;
  wire T20820;
  wire T20821;
  wire T20822;
  wire[46:0] T20823;
  wire[46:0] T20824;
  wire[46:0] T20825;
  wire[46:0] twiddle4_1_280_imag;
  wire[46:0] T20826;
  wire[46:0] T20827;
  wire[46:0] T20828;
  wire[46:0] T20829;
  wire[46:0] twiddle4_1_281_imag;
  wire[46:0] T20830;
  wire[46:0] T20831;
  wire[46:0] T20832;
  wire[46:0] T20833;
  wire T20834;
  wire[46:0] T20835;
  wire[46:0] twiddle4_1_282_imag;
  wire[46:0] T20836;
  wire[46:0] T20837;
  wire[46:0] T20838;
  wire[46:0] T20839;
  wire[46:0] twiddle4_1_283_imag;
  wire[46:0] T20840;
  wire[46:0] T20841;
  wire[46:0] T20842;
  wire[46:0] T20843;
  wire T20844;
  wire T20845;
  wire[46:0] T20846;
  wire[46:0] T20847;
  wire[46:0] twiddle4_1_284_imag;
  wire[46:0] T20848;
  wire[46:0] T20849;
  wire[46:0] T20850;
  wire[46:0] T20851;
  wire[46:0] twiddle4_1_285_imag;
  wire[46:0] T20852;
  wire[46:0] T20853;
  wire[46:0] T20854;
  wire[46:0] T20855;
  wire T20856;
  wire[46:0] T20857;
  wire[46:0] twiddle4_1_286_imag;
  wire[46:0] T20858;
  wire[46:0] T20859;
  wire[46:0] T20860;
  wire[46:0] T20861;
  wire[46:0] twiddle4_1_287_imag;
  wire[46:0] T20862;
  wire[46:0] T20863;
  wire[46:0] T20864;
  wire[46:0] T20865;
  wire T20866;
  wire T20867;
  wire T20868;
  wire T20869;
  wire T20870;
  wire[46:0] T20871;
  wire[46:0] T20872;
  wire[46:0] T20873;
  wire[46:0] T20874;
  wire[46:0] T20875;
  wire[46:0] twiddle4_1_288_imag;
  wire[46:0] T20876;
  wire[46:0] T20877;
  wire[46:0] T20878;
  wire[46:0] T20879;
  wire[46:0] twiddle4_1_289_imag;
  wire[46:0] T20880;
  wire[46:0] T20881;
  wire[46:0] T20882;
  wire[46:0] T20883;
  wire T20884;
  wire[46:0] T20885;
  wire[46:0] twiddle4_1_290_imag;
  wire[46:0] T20886;
  wire[46:0] T20887;
  wire[46:0] T20888;
  wire[46:0] T20889;
  wire[46:0] twiddle4_1_291_imag;
  wire[46:0] T20890;
  wire[46:0] T20891;
  wire[46:0] T20892;
  wire[46:0] T20893;
  wire T20894;
  wire T20895;
  wire[46:0] T20896;
  wire[46:0] T20897;
  wire[46:0] twiddle4_1_292_imag;
  wire[46:0] T20898;
  wire[46:0] T20899;
  wire[46:0] T20900;
  wire[46:0] T20901;
  wire[46:0] twiddle4_1_293_imag;
  wire[46:0] T20902;
  wire[46:0] T20903;
  wire[46:0] T20904;
  wire[46:0] T20905;
  wire T20906;
  wire[46:0] T20907;
  wire[46:0] twiddle4_1_294_imag;
  wire[46:0] T20908;
  wire[46:0] T20909;
  wire[46:0] T20910;
  wire[46:0] T20911;
  wire[46:0] twiddle4_1_295_imag;
  wire[46:0] T20912;
  wire[46:0] T20913;
  wire[46:0] T20914;
  wire[46:0] T20915;
  wire T20916;
  wire T20917;
  wire T20918;
  wire[46:0] T20919;
  wire[46:0] T20920;
  wire[46:0] T20921;
  wire[46:0] twiddle4_1_296_imag;
  wire[46:0] T20922;
  wire[46:0] T20923;
  wire[46:0] T20924;
  wire[46:0] T20925;
  wire[46:0] twiddle4_1_297_imag;
  wire[46:0] T20926;
  wire[46:0] T20927;
  wire[46:0] T20928;
  wire[46:0] T20929;
  wire T20930;
  wire[46:0] T20931;
  wire[46:0] twiddle4_1_298_imag;
  wire[46:0] T20932;
  wire[46:0] T20933;
  wire[46:0] T20934;
  wire[46:0] T20935;
  wire[46:0] twiddle4_1_299_imag;
  wire[46:0] T20936;
  wire[46:0] T20937;
  wire[46:0] T20938;
  wire[46:0] T20939;
  wire T20940;
  wire T20941;
  wire[46:0] T20942;
  wire[46:0] T20943;
  wire[46:0] twiddle4_1_300_imag;
  wire[46:0] T20944;
  wire[46:0] T20945;
  wire[46:0] T20946;
  wire[46:0] T20947;
  wire[46:0] twiddle4_1_301_imag;
  wire[46:0] T20948;
  wire[46:0] T20949;
  wire[46:0] T20950;
  wire[46:0] T20951;
  wire T20952;
  wire[46:0] T20953;
  wire[46:0] twiddle4_1_302_imag;
  wire[46:0] T20954;
  wire[46:0] T20955;
  wire[46:0] T20956;
  wire[46:0] T20957;
  wire[46:0] twiddle4_1_303_imag;
  wire[46:0] T20958;
  wire[46:0] T20959;
  wire[46:0] T20960;
  wire[46:0] T20961;
  wire T20962;
  wire T20963;
  wire T20964;
  wire T20965;
  wire[46:0] T20966;
  wire[46:0] T20967;
  wire[46:0] T20968;
  wire[46:0] T20969;
  wire[46:0] twiddle4_1_304_imag;
  wire[46:0] T20970;
  wire[46:0] T20971;
  wire[46:0] T20972;
  wire[46:0] T20973;
  wire[46:0] twiddle4_1_305_imag;
  wire[46:0] T20974;
  wire[46:0] T20975;
  wire[46:0] T20976;
  wire[46:0] T20977;
  wire T20978;
  wire[46:0] T20979;
  wire[46:0] twiddle4_1_306_imag;
  wire[46:0] T20980;
  wire[46:0] T20981;
  wire[46:0] T20982;
  wire[46:0] T20983;
  wire[46:0] twiddle4_1_307_imag;
  wire[46:0] T20984;
  wire[46:0] T20985;
  wire[46:0] T20986;
  wire[46:0] T20987;
  wire T20988;
  wire T20989;
  wire[46:0] T20990;
  wire[46:0] T20991;
  wire[46:0] twiddle4_1_308_imag;
  wire[46:0] T20992;
  wire[46:0] T20993;
  wire[46:0] T20994;
  wire[46:0] T20995;
  wire[46:0] twiddle4_1_309_imag;
  wire[46:0] T20996;
  wire[46:0] T20997;
  wire[46:0] T20998;
  wire[46:0] T20999;
  wire T21000;
  wire[46:0] T21001;
  wire[46:0] twiddle4_1_310_imag;
  wire[46:0] T21002;
  wire[46:0] T21003;
  wire[46:0] T21004;
  wire[46:0] T21005;
  wire[46:0] twiddle4_1_311_imag;
  wire[46:0] T21006;
  wire[46:0] T21007;
  wire[46:0] T21008;
  wire[46:0] T21009;
  wire T21010;
  wire T21011;
  wire T21012;
  wire[46:0] T21013;
  wire[46:0] T21014;
  wire[46:0] T21015;
  wire[46:0] twiddle4_1_312_imag;
  wire[46:0] T21016;
  wire[46:0] T21017;
  wire[46:0] T21018;
  wire[46:0] T21019;
  wire[46:0] twiddle4_1_313_imag;
  wire[46:0] T21020;
  wire[46:0] T21021;
  wire[46:0] T21022;
  wire[46:0] T21023;
  wire T21024;
  wire[46:0] T21025;
  wire[46:0] twiddle4_1_314_imag;
  wire[46:0] T21026;
  wire[46:0] T21027;
  wire[46:0] T21028;
  wire[46:0] T21029;
  wire[46:0] twiddle4_1_315_imag;
  wire[46:0] T21030;
  wire[46:0] T21031;
  wire[46:0] T21032;
  wire[46:0] T21033;
  wire T21034;
  wire T21035;
  wire[46:0] T21036;
  wire[46:0] T21037;
  wire[46:0] twiddle4_1_316_imag;
  wire[46:0] T21038;
  wire[46:0] T21039;
  wire[46:0] T21040;
  wire[46:0] T21041;
  wire[46:0] twiddle4_1_317_imag;
  wire[46:0] T21042;
  wire[46:0] T21043;
  wire[46:0] T21044;
  wire[46:0] T21045;
  wire T21046;
  wire[46:0] T21047;
  wire[46:0] twiddle4_1_318_imag;
  wire[46:0] T21048;
  wire[46:0] T21049;
  wire[46:0] T21050;
  wire[46:0] T21051;
  wire[46:0] twiddle4_1_319_imag;
  wire[46:0] T21052;
  wire[46:0] T21053;
  wire[46:0] T21054;
  wire[46:0] T21055;
  wire T21056;
  wire T21057;
  wire T21058;
  wire T21059;
  wire T21060;
  wire T21061;
  wire[46:0] T21062;
  wire[46:0] T21063;
  wire[46:0] T21064;
  wire[46:0] T21065;
  wire[46:0] T21066;
  wire[46:0] T21067;
  wire[46:0] twiddle4_1_320_imag;
  wire[46:0] T21068;
  wire[46:0] T21069;
  wire[46:0] T21070;
  wire[46:0] T21071;
  wire[46:0] twiddle4_1_321_imag;
  wire[46:0] T21072;
  wire[46:0] T21073;
  wire[46:0] T21074;
  wire[46:0] T21075;
  wire T21076;
  wire[46:0] T21077;
  wire[46:0] twiddle4_1_322_imag;
  wire[46:0] T21078;
  wire[46:0] T21079;
  wire[46:0] T21080;
  wire[46:0] T21081;
  wire[46:0] twiddle4_1_323_imag;
  wire[46:0] T21082;
  wire[46:0] T21083;
  wire[46:0] T21084;
  wire[46:0] T21085;
  wire T21086;
  wire T21087;
  wire[46:0] T21088;
  wire[46:0] T21089;
  wire[46:0] twiddle4_1_324_imag;
  wire[46:0] T21090;
  wire[46:0] T21091;
  wire[46:0] T21092;
  wire[46:0] T21093;
  wire[46:0] twiddle4_1_325_imag;
  wire[46:0] T21094;
  wire[46:0] T21095;
  wire[46:0] T21096;
  wire[46:0] T21097;
  wire T21098;
  wire[46:0] T21099;
  wire[46:0] twiddle4_1_326_imag;
  wire[46:0] T21100;
  wire[46:0] T21101;
  wire[46:0] T21102;
  wire[46:0] T21103;
  wire[46:0] twiddle4_1_327_imag;
  wire[46:0] T21104;
  wire[46:0] T21105;
  wire[46:0] T21106;
  wire[46:0] T21107;
  wire T21108;
  wire T21109;
  wire T21110;
  wire[46:0] T21111;
  wire[46:0] T21112;
  wire[46:0] T21113;
  wire[46:0] twiddle4_1_328_imag;
  wire[46:0] T21114;
  wire[46:0] T21115;
  wire[46:0] T21116;
  wire[46:0] T21117;
  wire[46:0] twiddle4_1_329_imag;
  wire[46:0] T21118;
  wire[46:0] T21119;
  wire[46:0] T21120;
  wire[46:0] T21121;
  wire T21122;
  wire[46:0] T21123;
  wire[46:0] twiddle4_1_330_imag;
  wire[46:0] T21124;
  wire[46:0] T21125;
  wire[46:0] T21126;
  wire[46:0] T21127;
  wire[46:0] twiddle4_1_331_imag;
  wire[46:0] T21128;
  wire[46:0] T21129;
  wire[46:0] T21130;
  wire[46:0] T21131;
  wire T21132;
  wire T21133;
  wire[46:0] T21134;
  wire[46:0] T21135;
  wire[46:0] twiddle4_1_332_imag;
  wire[46:0] T21136;
  wire[46:0] T21137;
  wire[46:0] T21138;
  wire[46:0] T21139;
  wire[46:0] twiddle4_1_333_imag;
  wire[46:0] T21140;
  wire[46:0] T21141;
  wire[46:0] T21142;
  wire[46:0] T21143;
  wire T21144;
  wire[46:0] T21145;
  wire[46:0] twiddle4_1_334_imag;
  wire[46:0] T21146;
  wire[46:0] T21147;
  wire[46:0] T21148;
  wire[46:0] T21149;
  wire[46:0] twiddle4_1_335_imag;
  wire[46:0] T21150;
  wire[46:0] T21151;
  wire[46:0] T21152;
  wire[46:0] T21153;
  wire T21154;
  wire T21155;
  wire T21156;
  wire T21157;
  wire[46:0] T21158;
  wire[46:0] T21159;
  wire[46:0] T21160;
  wire[46:0] T21161;
  wire[46:0] twiddle4_1_336_imag;
  wire[46:0] T21162;
  wire[46:0] T21163;
  wire[46:0] T21164;
  wire[46:0] T21165;
  wire[46:0] twiddle4_1_337_imag;
  wire[46:0] T21166;
  wire[46:0] T21167;
  wire[46:0] T21168;
  wire[46:0] T21169;
  wire T21170;
  wire[46:0] T21171;
  wire[46:0] twiddle4_1_338_imag;
  wire[46:0] T21172;
  wire[46:0] T21173;
  wire[46:0] T21174;
  wire[46:0] T21175;
  wire[46:0] twiddle4_1_339_imag;
  wire[46:0] T21176;
  wire[46:0] T21177;
  wire[46:0] T21178;
  wire[46:0] T21179;
  wire T21180;
  wire T21181;
  wire[46:0] T21182;
  wire[46:0] T21183;
  wire[46:0] twiddle4_1_340_imag;
  wire[46:0] T21184;
  wire[46:0] T21185;
  wire[46:0] T21186;
  wire[46:0] T21187;
  wire[46:0] twiddle4_1_341_imag;
  wire[46:0] T21188;
  wire[46:0] T21189;
  wire[46:0] T21190;
  wire[46:0] T21191;
  wire T21192;
  wire[46:0] T21193;
  wire[46:0] twiddle4_1_342_imag;
  wire[46:0] T21194;
  wire[46:0] T21195;
  wire[46:0] T21196;
  wire[45:0] T21197;
  wire[45:0] T21198;
  wire T21199;
  wire[46:0] twiddle4_1_343_imag;
  wire[46:0] T21200;
  wire[46:0] T21201;
  wire[46:0] T21202;
  wire[45:0] T21203;
  wire[45:0] T21204;
  wire T21205;
  wire T21206;
  wire T21207;
  wire T21208;
  wire[46:0] T21209;
  wire[46:0] T21210;
  wire[46:0] T21211;
  wire[46:0] twiddle4_1_344_imag;
  wire[46:0] T21212;
  wire[46:0] T21213;
  wire[46:0] T21214;
  wire[45:0] T21215;
  wire[45:0] T21216;
  wire T21217;
  wire[46:0] twiddle4_1_345_imag;
  wire[46:0] T21218;
  wire[46:0] T21219;
  wire[46:0] T21220;
  wire[45:0] T21221;
  wire[45:0] T21222;
  wire T21223;
  wire T21224;
  wire[46:0] T21225;
  wire[46:0] twiddle4_1_346_imag;
  wire[46:0] T21226;
  wire[46:0] T21227;
  wire[46:0] T21228;
  wire[45:0] T21229;
  wire[45:0] T21230;
  wire T21231;
  wire[46:0] twiddle4_1_347_imag;
  wire[46:0] T21232;
  wire[46:0] T21233;
  wire[46:0] T21234;
  wire[45:0] T21235;
  wire[45:0] T21236;
  wire T21237;
  wire T21238;
  wire T21239;
  wire[46:0] T21240;
  wire[46:0] T21241;
  wire[46:0] twiddle4_1_348_imag;
  wire[46:0] T21242;
  wire[46:0] T21243;
  wire[46:0] T21244;
  wire[45:0] T21245;
  wire[45:0] T21246;
  wire T21247;
  wire[46:0] twiddle4_1_349_imag;
  wire[46:0] T21248;
  wire[46:0] T21249;
  wire[46:0] T21250;
  wire[45:0] T21251;
  wire[45:0] T21252;
  wire T21253;
  wire T21254;
  wire[46:0] T21255;
  wire[46:0] twiddle4_1_350_imag;
  wire[46:0] T21256;
  wire[46:0] T21257;
  wire[46:0] T21258;
  wire[45:0] T21259;
  wire[45:0] T21260;
  wire T21261;
  wire[46:0] twiddle4_1_351_imag;
  wire[46:0] T21262;
  wire[46:0] T21263;
  wire[46:0] T21264;
  wire[45:0] T21265;
  wire[45:0] T21266;
  wire T21267;
  wire T21268;
  wire T21269;
  wire T21270;
  wire T21271;
  wire T21272;
  wire[46:0] T21273;
  wire[46:0] T21274;
  wire[46:0] T21275;
  wire[46:0] T21276;
  wire[46:0] T21277;
  wire[46:0] twiddle4_1_352_imag;
  wire[46:0] T21278;
  wire[46:0] T21279;
  wire[46:0] T21280;
  wire[45:0] T21281;
  wire[45:0] T21282;
  wire T21283;
  wire[46:0] twiddle4_1_353_imag;
  wire[46:0] T21284;
  wire[46:0] T21285;
  wire[46:0] T21286;
  wire[45:0] T21287;
  wire[45:0] T21288;
  wire T21289;
  wire T21290;
  wire[46:0] T21291;
  wire[46:0] twiddle4_1_354_imag;
  wire[46:0] T21292;
  wire[46:0] T21293;
  wire[46:0] T21294;
  wire[45:0] T21295;
  wire[45:0] T21296;
  wire T21297;
  wire[46:0] twiddle4_1_355_imag;
  wire[46:0] T21298;
  wire[46:0] T21299;
  wire[46:0] T21300;
  wire[45:0] T21301;
  wire[45:0] T21302;
  wire T21303;
  wire T21304;
  wire T21305;
  wire[46:0] T21306;
  wire[46:0] T21307;
  wire[46:0] twiddle4_1_356_imag;
  wire[46:0] T21308;
  wire[46:0] T21309;
  wire[46:0] T21310;
  wire[45:0] T21311;
  wire[45:0] T21312;
  wire T21313;
  wire[46:0] twiddle4_1_357_imag;
  wire[46:0] T21314;
  wire[46:0] T21315;
  wire[46:0] T21316;
  wire[45:0] T21317;
  wire[45:0] T21318;
  wire T21319;
  wire T21320;
  wire[46:0] T21321;
  wire[46:0] twiddle4_1_358_imag;
  wire[46:0] T21322;
  wire[46:0] T21323;
  wire[46:0] T21324;
  wire[45:0] T21325;
  wire[45:0] T21326;
  wire T21327;
  wire[46:0] twiddle4_1_359_imag;
  wire[46:0] T21328;
  wire[46:0] T21329;
  wire[46:0] T21330;
  wire[45:0] T21331;
  wire[45:0] T21332;
  wire T21333;
  wire T21334;
  wire T21335;
  wire T21336;
  wire[46:0] T21337;
  wire[46:0] T21338;
  wire[46:0] T21339;
  wire[46:0] twiddle4_1_360_imag;
  wire[46:0] T21340;
  wire[46:0] T21341;
  wire[46:0] T21342;
  wire[45:0] T21343;
  wire[45:0] T21344;
  wire T21345;
  wire[46:0] twiddle4_1_361_imag;
  wire[46:0] T21346;
  wire[46:0] T21347;
  wire[46:0] T21348;
  wire[45:0] T21349;
  wire[45:0] T21350;
  wire T21351;
  wire T21352;
  wire[46:0] T21353;
  wire[46:0] twiddle4_1_362_imag;
  wire[46:0] T21354;
  wire[46:0] T21355;
  wire[46:0] T21356;
  wire[45:0] T21357;
  wire[45:0] T21358;
  wire T21359;
  wire[46:0] twiddle4_1_363_imag;
  wire[46:0] T21360;
  wire[46:0] T21361;
  wire[46:0] T21362;
  wire[45:0] T21363;
  wire[45:0] T21364;
  wire T21365;
  wire T21366;
  wire T21367;
  wire[46:0] T21368;
  wire[46:0] T21369;
  wire[46:0] twiddle4_1_364_imag;
  wire[46:0] T21370;
  wire[46:0] T21371;
  wire[46:0] T21372;
  wire[45:0] T21373;
  wire[45:0] T21374;
  wire T21375;
  wire[46:0] twiddle4_1_365_imag;
  wire[46:0] T21376;
  wire[46:0] T21377;
  wire[46:0] T21378;
  wire[45:0] T21379;
  wire[45:0] T21380;
  wire T21381;
  wire T21382;
  wire[46:0] T21383;
  wire[46:0] twiddle4_1_366_imag;
  wire[46:0] T21384;
  wire[46:0] T21385;
  wire[46:0] T21386;
  wire[45:0] T21387;
  wire[45:0] T21388;
  wire T21389;
  wire[46:0] twiddle4_1_367_imag;
  wire[46:0] T21390;
  wire[46:0] T21391;
  wire[46:0] T21392;
  wire[45:0] T21393;
  wire[45:0] T21394;
  wire T21395;
  wire T21396;
  wire T21397;
  wire T21398;
  wire T21399;
  wire[46:0] T21400;
  wire[46:0] T21401;
  wire[46:0] T21402;
  wire[46:0] T21403;
  wire[46:0] twiddle4_1_368_imag;
  wire[46:0] T21404;
  wire[46:0] T21405;
  wire[46:0] T21406;
  wire[45:0] T21407;
  wire[45:0] T21408;
  wire T21409;
  wire[46:0] twiddle4_1_369_imag;
  wire[46:0] T21410;
  wire[46:0] T21411;
  wire[46:0] T21412;
  wire[45:0] T21413;
  wire[45:0] T21414;
  wire T21415;
  wire T21416;
  wire[46:0] T21417;
  wire[46:0] twiddle4_1_370_imag;
  wire[46:0] T21418;
  wire[46:0] T21419;
  wire[46:0] T21420;
  wire[45:0] T21421;
  wire[45:0] T21422;
  wire T21423;
  wire[46:0] twiddle4_1_371_imag;
  wire[46:0] T21424;
  wire[46:0] T21425;
  wire[46:0] T21426;
  wire[45:0] T21427;
  wire[45:0] T21428;
  wire T21429;
  wire T21430;
  wire T21431;
  wire[46:0] T21432;
  wire[46:0] T21433;
  wire[46:0] twiddle4_1_372_imag;
  wire[46:0] T21434;
  wire[46:0] T21435;
  wire[46:0] T21436;
  wire[45:0] T21437;
  wire[45:0] T21438;
  wire T21439;
  wire[46:0] twiddle4_1_373_imag;
  wire[46:0] T21440;
  wire[46:0] T21441;
  wire[46:0] T21442;
  wire[45:0] T21443;
  wire[45:0] T21444;
  wire T21445;
  wire T21446;
  wire[46:0] T21447;
  wire[46:0] twiddle4_1_374_imag;
  wire[46:0] T21448;
  wire[46:0] T21449;
  wire[46:0] T21450;
  wire[45:0] T21451;
  wire[45:0] T21452;
  wire T21453;
  wire[46:0] twiddle4_1_375_imag;
  wire[46:0] T21454;
  wire[46:0] T21455;
  wire[46:0] T21456;
  wire[45:0] T21457;
  wire[45:0] T21458;
  wire T21459;
  wire T21460;
  wire T21461;
  wire T21462;
  wire[46:0] T21463;
  wire[46:0] T21464;
  wire[46:0] T21465;
  wire[46:0] twiddle4_1_376_imag;
  wire[46:0] T21466;
  wire[46:0] T21467;
  wire[46:0] T21468;
  wire[45:0] T21469;
  wire[45:0] T21470;
  wire T21471;
  wire[46:0] twiddle4_1_377_imag;
  wire[46:0] T21472;
  wire[46:0] T21473;
  wire[46:0] T21474;
  wire[45:0] T21475;
  wire[45:0] T21476;
  wire T21477;
  wire T21478;
  wire[46:0] T21479;
  wire[46:0] twiddle4_1_378_imag;
  wire[46:0] T21480;
  wire[46:0] T21481;
  wire[46:0] T21482;
  wire[45:0] T21483;
  wire[45:0] T21484;
  wire T21485;
  wire[46:0] twiddle4_1_379_imag;
  wire[46:0] T21486;
  wire[46:0] T21487;
  wire[46:0] T21488;
  wire[45:0] T21489;
  wire[45:0] T21490;
  wire T21491;
  wire T21492;
  wire T21493;
  wire[46:0] T21494;
  wire[46:0] T21495;
  wire[46:0] twiddle4_1_380_imag;
  wire[46:0] T21496;
  wire[46:0] T21497;
  wire[46:0] T21498;
  wire[45:0] T21499;
  wire[45:0] T21500;
  wire T21501;
  wire[46:0] twiddle4_1_381_imag;
  wire[46:0] T21502;
  wire[46:0] T21503;
  wire[46:0] T21504;
  wire[45:0] T21505;
  wire[45:0] T21506;
  wire T21507;
  wire T21508;
  wire[46:0] T21509;
  wire[46:0] twiddle4_1_382_imag;
  wire[46:0] T21510;
  wire[46:0] T21511;
  wire[46:0] T21512;
  wire[45:0] T21513;
  wire[45:0] T21514;
  wire T21515;
  wire[46:0] twiddle4_1_383_imag;
  wire[46:0] T21516;
  wire[46:0] T21517;
  wire[46:0] T21518;
  wire[45:0] T21519;
  wire[45:0] T21520;
  wire T21521;
  wire T21522;
  wire T21523;
  wire T21524;
  wire T21525;
  wire T21526;
  wire T21527;
  wire T21528;
  wire[46:0] T21529;
  wire[46:0] T21530;
  wire[46:0] T21531;
  wire[46:0] T21532;
  wire[46:0] T21533;
  wire[46:0] T21534;
  wire[46:0] T21535;
  wire[46:0] twiddle4_1_384_imag;
  wire[46:0] T21536;
  wire[46:0] T21537;
  wire[46:0] T21538;
  wire[45:0] T21539;
  wire[45:0] T21540;
  wire T21541;
  wire[46:0] twiddle4_1_385_imag;
  wire[46:0] T21542;
  wire[46:0] T21543;
  wire[46:0] T21544;
  wire[45:0] T21545;
  wire[45:0] T21546;
  wire T21547;
  wire T21548;
  wire[46:0] T21549;
  wire[46:0] twiddle4_1_386_imag;
  wire[46:0] T21550;
  wire[46:0] T21551;
  wire[46:0] T21552;
  wire[45:0] T21553;
  wire[45:0] T21554;
  wire T21555;
  wire[46:0] twiddle4_1_387_imag;
  wire[46:0] T21556;
  wire[46:0] T21557;
  wire[46:0] T21558;
  wire[45:0] T21559;
  wire[45:0] T21560;
  wire T21561;
  wire T21562;
  wire T21563;
  wire[46:0] T21564;
  wire[46:0] T21565;
  wire[46:0] twiddle4_1_388_imag;
  wire[46:0] T21566;
  wire[46:0] T21567;
  wire[46:0] T21568;
  wire[45:0] T21569;
  wire[45:0] T21570;
  wire T21571;
  wire[46:0] twiddle4_1_389_imag;
  wire[46:0] T21572;
  wire[46:0] T21573;
  wire[46:0] T21574;
  wire[45:0] T21575;
  wire[45:0] T21576;
  wire T21577;
  wire T21578;
  wire[46:0] T21579;
  wire[46:0] twiddle4_1_390_imag;
  wire[46:0] T21580;
  wire[46:0] T21581;
  wire[46:0] T21582;
  wire[45:0] T21583;
  wire[45:0] T21584;
  wire T21585;
  wire[46:0] twiddle4_1_391_imag;
  wire[46:0] T21586;
  wire[46:0] T21587;
  wire[46:0] T21588;
  wire[45:0] T21589;
  wire[45:0] T21590;
  wire T21591;
  wire T21592;
  wire T21593;
  wire T21594;
  wire[46:0] T21595;
  wire[46:0] T21596;
  wire[46:0] T21597;
  wire[46:0] twiddle4_1_392_imag;
  wire[46:0] T21598;
  wire[46:0] T21599;
  wire[46:0] T21600;
  wire[45:0] T21601;
  wire[45:0] T21602;
  wire T21603;
  wire[46:0] twiddle4_1_393_imag;
  wire[46:0] T21604;
  wire[46:0] T21605;
  wire[46:0] T21606;
  wire[45:0] T21607;
  wire[45:0] T21608;
  wire T21609;
  wire T21610;
  wire[46:0] T21611;
  wire[46:0] twiddle4_1_394_imag;
  wire[46:0] T21612;
  wire[46:0] T21613;
  wire[46:0] T21614;
  wire[45:0] T21615;
  wire[45:0] T21616;
  wire T21617;
  wire[46:0] twiddle4_1_395_imag;
  wire[46:0] T21618;
  wire[46:0] T21619;
  wire[46:0] T21620;
  wire[45:0] T21621;
  wire[45:0] T21622;
  wire T21623;
  wire T21624;
  wire T21625;
  wire[46:0] T21626;
  wire[46:0] T21627;
  wire[46:0] twiddle4_1_396_imag;
  wire[46:0] T21628;
  wire[46:0] T21629;
  wire[46:0] T21630;
  wire[45:0] T21631;
  wire[45:0] T21632;
  wire T21633;
  wire[46:0] twiddle4_1_397_imag;
  wire[46:0] T21634;
  wire[46:0] T21635;
  wire[46:0] T21636;
  wire[45:0] T21637;
  wire[45:0] T21638;
  wire T21639;
  wire T21640;
  wire[46:0] T21641;
  wire[46:0] twiddle4_1_398_imag;
  wire[46:0] T21642;
  wire[46:0] T21643;
  wire[46:0] T21644;
  wire[45:0] T21645;
  wire[45:0] T21646;
  wire T21647;
  wire[46:0] twiddle4_1_399_imag;
  wire[46:0] T21648;
  wire[46:0] T21649;
  wire[46:0] T21650;
  wire[45:0] T21651;
  wire[45:0] T21652;
  wire T21653;
  wire T21654;
  wire T21655;
  wire T21656;
  wire T21657;
  wire[46:0] T21658;
  wire[46:0] T21659;
  wire[46:0] T21660;
  wire[46:0] T21661;
  wire[46:0] twiddle4_1_400_imag;
  wire[46:0] T21662;
  wire[46:0] T21663;
  wire[46:0] T21664;
  wire[45:0] T21665;
  wire[45:0] T21666;
  wire T21667;
  wire[46:0] twiddle4_1_401_imag;
  wire[46:0] T21668;
  wire[46:0] T21669;
  wire[46:0] T21670;
  wire[45:0] T21671;
  wire[45:0] T21672;
  wire T21673;
  wire T21674;
  wire[46:0] T21675;
  wire[46:0] twiddle4_1_402_imag;
  wire[46:0] T21676;
  wire[46:0] T21677;
  wire[46:0] T21678;
  wire[45:0] T21679;
  wire[45:0] T21680;
  wire T21681;
  wire[46:0] twiddle4_1_403_imag;
  wire[46:0] T21682;
  wire[46:0] T21683;
  wire[46:0] T21684;
  wire[45:0] T21685;
  wire[45:0] T21686;
  wire T21687;
  wire T21688;
  wire T21689;
  wire[46:0] T21690;
  wire[46:0] T21691;
  wire[46:0] twiddle4_1_404_imag;
  wire[46:0] T21692;
  wire[46:0] T21693;
  wire[46:0] T21694;
  wire[45:0] T21695;
  wire[45:0] T21696;
  wire T21697;
  wire[46:0] twiddle4_1_405_imag;
  wire[46:0] T21698;
  wire[46:0] T21699;
  wire[46:0] T21700;
  wire[45:0] T21701;
  wire[45:0] T21702;
  wire T21703;
  wire T21704;
  wire[46:0] T21705;
  wire[46:0] twiddle4_1_406_imag;
  wire[46:0] T21706;
  wire[46:0] T21707;
  wire[46:0] T21708;
  wire[45:0] T21709;
  wire[45:0] T21710;
  wire T21711;
  wire[46:0] twiddle4_1_407_imag;
  wire[46:0] T21712;
  wire[46:0] T21713;
  wire[46:0] T21714;
  wire[45:0] T21715;
  wire[45:0] T21716;
  wire T21717;
  wire T21718;
  wire T21719;
  wire T21720;
  wire[46:0] T21721;
  wire[46:0] T21722;
  wire[46:0] T21723;
  wire[46:0] twiddle4_1_408_imag;
  wire[46:0] T21724;
  wire[46:0] T21725;
  wire[46:0] T21726;
  wire[45:0] T21727;
  wire[45:0] T21728;
  wire T21729;
  wire[46:0] twiddle4_1_409_imag;
  wire[46:0] T21730;
  wire[46:0] T21731;
  wire[46:0] T21732;
  wire[45:0] T21733;
  wire[45:0] T21734;
  wire T21735;
  wire T21736;
  wire[46:0] T21737;
  wire[46:0] twiddle4_1_410_imag;
  wire[46:0] T21738;
  wire[46:0] T21739;
  wire[46:0] T21740;
  wire[45:0] T21741;
  wire[45:0] T21742;
  wire T21743;
  wire[46:0] twiddle4_1_411_imag;
  wire[46:0] T21744;
  wire[46:0] T21745;
  wire[46:0] T21746;
  wire[45:0] T21747;
  wire[45:0] T21748;
  wire T21749;
  wire T21750;
  wire T21751;
  wire[46:0] T21752;
  wire[46:0] T21753;
  wire[46:0] twiddle4_1_412_imag;
  wire[46:0] T21754;
  wire[46:0] T21755;
  wire[46:0] T21756;
  wire[45:0] T21757;
  wire[45:0] T21758;
  wire T21759;
  wire[46:0] twiddle4_1_413_imag;
  wire[46:0] T21760;
  wire[46:0] T21761;
  wire[46:0] T21762;
  wire[45:0] T21763;
  wire[45:0] T21764;
  wire T21765;
  wire T21766;
  wire[46:0] T21767;
  wire[46:0] twiddle4_1_414_imag;
  wire[46:0] T21768;
  wire[46:0] T21769;
  wire[46:0] T21770;
  wire[45:0] T21771;
  wire[45:0] T21772;
  wire T21773;
  wire[46:0] twiddle4_1_415_imag;
  wire[46:0] T21774;
  wire[46:0] T21775;
  wire[46:0] T21776;
  wire[45:0] T21777;
  wire[45:0] T21778;
  wire T21779;
  wire T21780;
  wire T21781;
  wire T21782;
  wire T21783;
  wire T21784;
  wire[46:0] T21785;
  wire[46:0] T21786;
  wire[46:0] T21787;
  wire[46:0] T21788;
  wire[46:0] T21789;
  wire[46:0] twiddle4_1_416_imag;
  wire[46:0] T21790;
  wire[46:0] T21791;
  wire[46:0] T21792;
  wire[45:0] T21793;
  wire[45:0] T21794;
  wire T21795;
  wire[46:0] twiddle4_1_417_imag;
  wire[46:0] T21796;
  wire[46:0] T21797;
  wire[46:0] T21798;
  wire[45:0] T21799;
  wire[45:0] T21800;
  wire T21801;
  wire T21802;
  wire[46:0] T21803;
  wire[46:0] twiddle4_1_418_imag;
  wire[46:0] T21804;
  wire[46:0] T21805;
  wire[46:0] T21806;
  wire[45:0] T21807;
  wire[45:0] T21808;
  wire T21809;
  wire[46:0] twiddle4_1_419_imag;
  wire[46:0] T21810;
  wire[46:0] T21811;
  wire[46:0] T21812;
  wire[45:0] T21813;
  wire[45:0] T21814;
  wire T21815;
  wire T21816;
  wire T21817;
  wire[46:0] T21818;
  wire[46:0] T21819;
  wire[46:0] twiddle4_1_420_imag;
  wire[46:0] T21820;
  wire[46:0] T21821;
  wire[46:0] T21822;
  wire[45:0] T21823;
  wire[45:0] T21824;
  wire T21825;
  wire[46:0] twiddle4_1_421_imag;
  wire[46:0] T21826;
  wire[46:0] T21827;
  wire[46:0] T21828;
  wire[45:0] T21829;
  wire[45:0] T21830;
  wire T21831;
  wire T21832;
  wire[46:0] T21833;
  wire[46:0] twiddle4_1_422_imag;
  wire[46:0] T21834;
  wire[46:0] T21835;
  wire[46:0] T21836;
  wire[45:0] T21837;
  wire[45:0] T21838;
  wire T21839;
  wire[46:0] twiddle4_1_423_imag;
  wire[46:0] T21840;
  wire[46:0] T21841;
  wire[46:0] T21842;
  wire[45:0] T21843;
  wire[45:0] T21844;
  wire T21845;
  wire T21846;
  wire T21847;
  wire T21848;
  wire[46:0] T21849;
  wire[46:0] T21850;
  wire[46:0] T21851;
  wire[46:0] twiddle4_1_424_imag;
  wire[46:0] T21852;
  wire[46:0] T21853;
  wire[46:0] T21854;
  wire[45:0] T21855;
  wire[45:0] T21856;
  wire T21857;
  wire[46:0] twiddle4_1_425_imag;
  wire[46:0] T21858;
  wire[46:0] T21859;
  wire[46:0] T21860;
  wire[45:0] T21861;
  wire[45:0] T21862;
  wire T21863;
  wire T21864;
  wire[46:0] T21865;
  wire[46:0] twiddle4_1_426_imag;
  wire[46:0] T21866;
  wire[46:0] T21867;
  wire[46:0] T21868;
  wire[45:0] T21869;
  wire[45:0] T21870;
  wire T21871;
  wire[46:0] twiddle4_1_427_imag;
  wire[46:0] T21872;
  wire[46:0] T21873;
  wire[46:0] T21874;
  wire[45:0] T21875;
  wire[45:0] T21876;
  wire T21877;
  wire T21878;
  wire T21879;
  wire[46:0] T21880;
  wire[46:0] T21881;
  wire[46:0] twiddle4_1_428_imag;
  wire[46:0] T21882;
  wire[46:0] T21883;
  wire[46:0] T21884;
  wire[45:0] T21885;
  wire[45:0] T21886;
  wire T21887;
  wire[46:0] twiddle4_1_429_imag;
  wire[46:0] T21888;
  wire[46:0] T21889;
  wire[46:0] T21890;
  wire[45:0] T21891;
  wire[45:0] T21892;
  wire T21893;
  wire T21894;
  wire[46:0] T21895;
  wire[46:0] twiddle4_1_430_imag;
  wire[46:0] T21896;
  wire[46:0] T21897;
  wire[46:0] T21898;
  wire[44:0] T21899;
  wire[44:0] T21900;
  wire[1:0] T21901;
  wire T21902;
  wire[46:0] twiddle4_1_431_imag;
  wire[46:0] T21903;
  wire[46:0] T21904;
  wire[46:0] T21905;
  wire[44:0] T21906;
  wire[44:0] T21907;
  wire[1:0] T21908;
  wire T21909;
  wire T21910;
  wire T21911;
  wire T21912;
  wire T21913;
  wire[46:0] T21914;
  wire[46:0] T21915;
  wire[46:0] T21916;
  wire[46:0] T21917;
  wire[46:0] twiddle4_1_432_imag;
  wire[46:0] T21918;
  wire[46:0] T21919;
  wire[46:0] T21920;
  wire[44:0] T21921;
  wire[44:0] T21922;
  wire[1:0] T21923;
  wire T21924;
  wire[46:0] twiddle4_1_433_imag;
  wire[46:0] T21925;
  wire[46:0] T21926;
  wire[46:0] T21927;
  wire[44:0] T21928;
  wire[44:0] T21929;
  wire[1:0] T21930;
  wire T21931;
  wire T21932;
  wire[46:0] T21933;
  wire[46:0] twiddle4_1_434_imag;
  wire[46:0] T21934;
  wire[46:0] T21935;
  wire[46:0] T21936;
  wire[44:0] T21937;
  wire[44:0] T21938;
  wire[1:0] T21939;
  wire T21940;
  wire[46:0] twiddle4_1_435_imag;
  wire[46:0] T21941;
  wire[46:0] T21942;
  wire[46:0] T21943;
  wire[44:0] T21944;
  wire[44:0] T21945;
  wire[1:0] T21946;
  wire T21947;
  wire T21948;
  wire T21949;
  wire[46:0] T21950;
  wire[46:0] T21951;
  wire[46:0] twiddle4_1_436_imag;
  wire[46:0] T21952;
  wire[46:0] T21953;
  wire[46:0] T21954;
  wire[44:0] T21955;
  wire[44:0] T21956;
  wire[1:0] T21957;
  wire T21958;
  wire[46:0] twiddle4_1_437_imag;
  wire[46:0] T21959;
  wire[46:0] T21960;
  wire[46:0] T21961;
  wire[44:0] T21962;
  wire[44:0] T21963;
  wire[1:0] T21964;
  wire T21965;
  wire T21966;
  wire[46:0] T21967;
  wire[46:0] twiddle4_1_438_imag;
  wire[46:0] T21968;
  wire[46:0] T21969;
  wire[46:0] T21970;
  wire[44:0] T21971;
  wire[44:0] T21972;
  wire[1:0] T21973;
  wire T21974;
  wire[46:0] twiddle4_1_439_imag;
  wire[46:0] T21975;
  wire[46:0] T21976;
  wire[46:0] T21977;
  wire[44:0] T21978;
  wire[44:0] T21979;
  wire[1:0] T21980;
  wire T21981;
  wire T21982;
  wire T21983;
  wire T21984;
  wire[46:0] T21985;
  wire[46:0] T21986;
  wire[46:0] T21987;
  wire[46:0] twiddle4_1_440_imag;
  wire[46:0] T21988;
  wire[46:0] T21989;
  wire[46:0] T21990;
  wire[44:0] T21991;
  wire[44:0] T21992;
  wire[1:0] T21993;
  wire T21994;
  wire[46:0] twiddle4_1_441_imag;
  wire[46:0] T21995;
  wire[46:0] T21996;
  wire[46:0] T21997;
  wire[44:0] T21998;
  wire[44:0] T21999;
  wire[1:0] T22000;
  wire T22001;
  wire T22002;
  wire[46:0] T22003;
  wire[46:0] twiddle4_1_442_imag;
  wire[46:0] T22004;
  wire[46:0] T22005;
  wire[46:0] T22006;
  wire[44:0] T22007;
  wire[44:0] T22008;
  wire[1:0] T22009;
  wire T22010;
  wire[46:0] twiddle4_1_443_imag;
  wire[46:0] T22011;
  wire[46:0] T22012;
  wire[46:0] T22013;
  wire[44:0] T22014;
  wire[44:0] T22015;
  wire[1:0] T22016;
  wire T22017;
  wire T22018;
  wire T22019;
  wire[46:0] T22020;
  wire[46:0] T22021;
  wire[46:0] twiddle4_1_444_imag;
  wire[46:0] T22022;
  wire[46:0] T22023;
  wire[46:0] T22024;
  wire[44:0] T22025;
  wire[44:0] T22026;
  wire[1:0] T22027;
  wire T22028;
  wire[46:0] twiddle4_1_445_imag;
  wire[46:0] T22029;
  wire[46:0] T22030;
  wire[46:0] T22031;
  wire[44:0] T22032;
  wire[44:0] T22033;
  wire[1:0] T22034;
  wire T22035;
  wire T22036;
  wire[46:0] T22037;
  wire[46:0] twiddle4_1_446_imag;
  wire[46:0] T22038;
  wire[46:0] T22039;
  wire[46:0] T22040;
  wire[44:0] T22041;
  wire[44:0] T22042;
  wire[1:0] T22043;
  wire T22044;
  wire[46:0] twiddle4_1_447_imag;
  wire[46:0] T22045;
  wire[46:0] T22046;
  wire[46:0] T22047;
  wire[44:0] T22048;
  wire[44:0] T22049;
  wire[1:0] T22050;
  wire T22051;
  wire T22052;
  wire T22053;
  wire T22054;
  wire T22055;
  wire T22056;
  wire T22057;
  wire[46:0] T22058;
  wire[46:0] T22059;
  wire[46:0] T22060;
  wire[46:0] T22061;
  wire[46:0] T22062;
  wire[46:0] T22063;
  wire[46:0] twiddle4_1_448_imag;
  wire[46:0] T22064;
  wire[46:0] T22065;
  wire[46:0] T22066;
  wire[44:0] T22067;
  wire[44:0] T22068;
  wire[1:0] T22069;
  wire T22070;
  wire[46:0] twiddle4_1_449_imag;
  wire[46:0] T22071;
  wire[46:0] T22072;
  wire[46:0] T22073;
  wire[44:0] T22074;
  wire[44:0] T22075;
  wire[1:0] T22076;
  wire T22077;
  wire T22078;
  wire[46:0] T22079;
  wire[46:0] twiddle4_1_450_imag;
  wire[46:0] T22080;
  wire[46:0] T22081;
  wire[46:0] T22082;
  wire[44:0] T22083;
  wire[44:0] T22084;
  wire[1:0] T22085;
  wire T22086;
  wire[46:0] twiddle4_1_451_imag;
  wire[46:0] T22087;
  wire[46:0] T22088;
  wire[46:0] T22089;
  wire[44:0] T22090;
  wire[44:0] T22091;
  wire[1:0] T22092;
  wire T22093;
  wire T22094;
  wire T22095;
  wire[46:0] T22096;
  wire[46:0] T22097;
  wire[46:0] twiddle4_1_452_imag;
  wire[46:0] T22098;
  wire[46:0] T22099;
  wire[46:0] T22100;
  wire[44:0] T22101;
  wire[44:0] T22102;
  wire[1:0] T22103;
  wire T22104;
  wire[46:0] twiddle4_1_453_imag;
  wire[46:0] T22105;
  wire[46:0] T22106;
  wire[46:0] T22107;
  wire[44:0] T22108;
  wire[44:0] T22109;
  wire[1:0] T22110;
  wire T22111;
  wire T22112;
  wire[46:0] T22113;
  wire[46:0] twiddle4_1_454_imag;
  wire[46:0] T22114;
  wire[46:0] T22115;
  wire[46:0] T22116;
  wire[44:0] T22117;
  wire[44:0] T22118;
  wire[1:0] T22119;
  wire T22120;
  wire[46:0] twiddle4_1_455_imag;
  wire[46:0] T22121;
  wire[46:0] T22122;
  wire[46:0] T22123;
  wire[44:0] T22124;
  wire[44:0] T22125;
  wire[1:0] T22126;
  wire T22127;
  wire T22128;
  wire T22129;
  wire T22130;
  wire[46:0] T22131;
  wire[46:0] T22132;
  wire[46:0] T22133;
  wire[46:0] twiddle4_1_456_imag;
  wire[46:0] T22134;
  wire[46:0] T22135;
  wire[46:0] T22136;
  wire[44:0] T22137;
  wire[44:0] T22138;
  wire[1:0] T22139;
  wire T22140;
  wire[46:0] twiddle4_1_457_imag;
  wire[46:0] T22141;
  wire[46:0] T22142;
  wire[46:0] T22143;
  wire[44:0] T22144;
  wire[44:0] T22145;
  wire[1:0] T22146;
  wire T22147;
  wire T22148;
  wire[46:0] T22149;
  wire[46:0] twiddle4_1_458_imag;
  wire[46:0] T22150;
  wire[46:0] T22151;
  wire[46:0] T22152;
  wire[44:0] T22153;
  wire[44:0] T22154;
  wire[1:0] T22155;
  wire T22156;
  wire[46:0] twiddle4_1_459_imag;
  wire[46:0] T22157;
  wire[46:0] T22158;
  wire[46:0] T22159;
  wire[44:0] T22160;
  wire[44:0] T22161;
  wire[1:0] T22162;
  wire T22163;
  wire T22164;
  wire T22165;
  wire[46:0] T22166;
  wire[46:0] T22167;
  wire[46:0] twiddle4_1_460_imag;
  wire[46:0] T22168;
  wire[46:0] T22169;
  wire[46:0] T22170;
  wire[44:0] T22171;
  wire[44:0] T22172;
  wire[1:0] T22173;
  wire T22174;
  wire[46:0] twiddle4_1_461_imag;
  wire[46:0] T22175;
  wire[46:0] T22176;
  wire[46:0] T22177;
  wire[44:0] T22178;
  wire[44:0] T22179;
  wire[1:0] T22180;
  wire T22181;
  wire T22182;
  wire[46:0] T22183;
  wire[46:0] twiddle4_1_462_imag;
  wire[46:0] T22184;
  wire[46:0] T22185;
  wire[46:0] T22186;
  wire[44:0] T22187;
  wire[44:0] T22188;
  wire[1:0] T22189;
  wire T22190;
  wire[46:0] twiddle4_1_463_imag;
  wire[46:0] T22191;
  wire[46:0] T22192;
  wire[46:0] T22193;
  wire[44:0] T22194;
  wire[44:0] T22195;
  wire[1:0] T22196;
  wire T22197;
  wire T22198;
  wire T22199;
  wire T22200;
  wire T22201;
  wire[46:0] T22202;
  wire[46:0] T22203;
  wire[46:0] T22204;
  wire[46:0] T22205;
  wire[46:0] twiddle4_1_464_imag;
  wire[46:0] T22206;
  wire[46:0] T22207;
  wire[46:0] T22208;
  wire[44:0] T22209;
  wire[44:0] T22210;
  wire[1:0] T22211;
  wire T22212;
  wire[46:0] twiddle4_1_465_imag;
  wire[46:0] T22213;
  wire[46:0] T22214;
  wire[46:0] T22215;
  wire[44:0] T22216;
  wire[44:0] T22217;
  wire[1:0] T22218;
  wire T22219;
  wire T22220;
  wire[46:0] T22221;
  wire[46:0] twiddle4_1_466_imag;
  wire[46:0] T22222;
  wire[46:0] T22223;
  wire[46:0] T22224;
  wire[44:0] T22225;
  wire[44:0] T22226;
  wire[1:0] T22227;
  wire T22228;
  wire[46:0] twiddle4_1_467_imag;
  wire[46:0] T22229;
  wire[46:0] T22230;
  wire[46:0] T22231;
  wire[44:0] T22232;
  wire[44:0] T22233;
  wire[1:0] T22234;
  wire T22235;
  wire T22236;
  wire T22237;
  wire[46:0] T22238;
  wire[46:0] T22239;
  wire[46:0] twiddle4_1_468_imag;
  wire[46:0] T22240;
  wire[46:0] T22241;
  wire[46:0] T22242;
  wire[44:0] T22243;
  wire[44:0] T22244;
  wire[1:0] T22245;
  wire T22246;
  wire[46:0] twiddle4_1_469_imag;
  wire[46:0] T22247;
  wire[46:0] T22248;
  wire[46:0] T22249;
  wire[44:0] T22250;
  wire[44:0] T22251;
  wire[1:0] T22252;
  wire T22253;
  wire T22254;
  wire[46:0] T22255;
  wire[46:0] twiddle4_1_470_imag;
  wire[46:0] T22256;
  wire[46:0] T22257;
  wire[46:0] T22258;
  wire[44:0] T22259;
  wire[44:0] T22260;
  wire[1:0] T22261;
  wire T22262;
  wire[46:0] twiddle4_1_471_imag;
  wire[46:0] T22263;
  wire[46:0] T22264;
  wire[46:0] T22265;
  wire[44:0] T22266;
  wire[44:0] T22267;
  wire[1:0] T22268;
  wire T22269;
  wire T22270;
  wire T22271;
  wire T22272;
  wire[46:0] T22273;
  wire[46:0] T22274;
  wire[46:0] T22275;
  wire[46:0] twiddle4_1_472_imag;
  wire[46:0] T22276;
  wire[46:0] T22277;
  wire[46:0] T22278;
  wire[43:0] T22279;
  wire[43:0] T22280;
  wire[2:0] T22281;
  wire T22282;
  wire[46:0] twiddle4_1_473_imag;
  wire[46:0] T22283;
  wire[46:0] T22284;
  wire[46:0] T22285;
  wire[43:0] T22286;
  wire[43:0] T22287;
  wire[2:0] T22288;
  wire T22289;
  wire T22290;
  wire[46:0] T22291;
  wire[46:0] twiddle4_1_474_imag;
  wire[46:0] T22292;
  wire[46:0] T22293;
  wire[46:0] T22294;
  wire[43:0] T22295;
  wire[43:0] T22296;
  wire[2:0] T22297;
  wire T22298;
  wire[46:0] twiddle4_1_475_imag;
  wire[46:0] T22299;
  wire[46:0] T22300;
  wire[46:0] T22301;
  wire[43:0] T22302;
  wire[43:0] T22303;
  wire[2:0] T22304;
  wire T22305;
  wire T22306;
  wire T22307;
  wire[46:0] T22308;
  wire[46:0] T22309;
  wire[46:0] twiddle4_1_476_imag;
  wire[46:0] T22310;
  wire[46:0] T22311;
  wire[46:0] T22312;
  wire[43:0] T22313;
  wire[43:0] T22314;
  wire[2:0] T22315;
  wire T22316;
  wire[46:0] twiddle4_1_477_imag;
  wire[46:0] T22317;
  wire[46:0] T22318;
  wire[46:0] T22319;
  wire[43:0] T22320;
  wire[43:0] T22321;
  wire[2:0] T22322;
  wire T22323;
  wire T22324;
  wire[46:0] T22325;
  wire[46:0] twiddle4_1_478_imag;
  wire[46:0] T22326;
  wire[46:0] T22327;
  wire[46:0] T22328;
  wire[43:0] T22329;
  wire[43:0] T22330;
  wire[2:0] T22331;
  wire T22332;
  wire[46:0] twiddle4_1_479_imag;
  wire[46:0] T22333;
  wire[46:0] T22334;
  wire[46:0] T22335;
  wire[43:0] T22336;
  wire[43:0] T22337;
  wire[2:0] T22338;
  wire T22339;
  wire T22340;
  wire T22341;
  wire T22342;
  wire T22343;
  wire T22344;
  wire[46:0] T22345;
  wire[46:0] T22346;
  wire[46:0] T22347;
  wire[46:0] T22348;
  wire[46:0] T22349;
  wire[46:0] twiddle4_1_480_imag;
  wire[46:0] T22350;
  wire[46:0] T22351;
  wire[46:0] T22352;
  wire[43:0] T22353;
  wire[43:0] T22354;
  wire[2:0] T22355;
  wire T22356;
  wire[46:0] twiddle4_1_481_imag;
  wire[46:0] T22357;
  wire[46:0] T22358;
  wire[46:0] T22359;
  wire[43:0] T22360;
  wire[43:0] T22361;
  wire[2:0] T22362;
  wire T22363;
  wire T22364;
  wire[46:0] T22365;
  wire[46:0] twiddle4_1_482_imag;
  wire[46:0] T22366;
  wire[46:0] T22367;
  wire[46:0] T22368;
  wire[43:0] T22369;
  wire[43:0] T22370;
  wire[2:0] T22371;
  wire T22372;
  wire[46:0] twiddle4_1_483_imag;
  wire[46:0] T22373;
  wire[46:0] T22374;
  wire[46:0] T22375;
  wire[43:0] T22376;
  wire[43:0] T22377;
  wire[2:0] T22378;
  wire T22379;
  wire T22380;
  wire T22381;
  wire[46:0] T22382;
  wire[46:0] T22383;
  wire[46:0] twiddle4_1_484_imag;
  wire[46:0] T22384;
  wire[46:0] T22385;
  wire[46:0] T22386;
  wire[43:0] T22387;
  wire[43:0] T22388;
  wire[2:0] T22389;
  wire T22390;
  wire[46:0] twiddle4_1_485_imag;
  wire[46:0] T22391;
  wire[46:0] T22392;
  wire[46:0] T22393;
  wire[43:0] T22394;
  wire[43:0] T22395;
  wire[2:0] T22396;
  wire T22397;
  wire T22398;
  wire[46:0] T22399;
  wire[46:0] twiddle4_1_486_imag;
  wire[46:0] T22400;
  wire[46:0] T22401;
  wire[46:0] T22402;
  wire[43:0] T22403;
  wire[43:0] T22404;
  wire[2:0] T22405;
  wire T22406;
  wire[46:0] twiddle4_1_487_imag;
  wire[46:0] T22407;
  wire[46:0] T22408;
  wire[46:0] T22409;
  wire[43:0] T22410;
  wire[43:0] T22411;
  wire[2:0] T22412;
  wire T22413;
  wire T22414;
  wire T22415;
  wire T22416;
  wire[46:0] T22417;
  wire[46:0] T22418;
  wire[46:0] T22419;
  wire[46:0] twiddle4_1_488_imag;
  wire[46:0] T22420;
  wire[46:0] T22421;
  wire[46:0] T22422;
  wire[43:0] T22423;
  wire[43:0] T22424;
  wire[2:0] T22425;
  wire T22426;
  wire[46:0] twiddle4_1_489_imag;
  wire[46:0] T22427;
  wire[46:0] T22428;
  wire[46:0] T22429;
  wire[43:0] T22430;
  wire[43:0] T22431;
  wire[2:0] T22432;
  wire T22433;
  wire T22434;
  wire[46:0] T22435;
  wire[46:0] twiddle4_1_490_imag;
  wire[46:0] T22436;
  wire[46:0] T22437;
  wire[46:0] T22438;
  wire[43:0] T22439;
  wire[43:0] T22440;
  wire[2:0] T22441;
  wire T22442;
  wire[46:0] twiddle4_1_491_imag;
  wire[46:0] T22443;
  wire[46:0] T22444;
  wire[46:0] T22445;
  wire[43:0] T22446;
  wire[43:0] T22447;
  wire[2:0] T22448;
  wire T22449;
  wire T22450;
  wire T22451;
  wire[46:0] T22452;
  wire[46:0] T22453;
  wire[46:0] twiddle4_1_492_imag;
  wire[46:0] T22454;
  wire[46:0] T22455;
  wire[46:0] T22456;
  wire[42:0] T22457;
  wire[42:0] T22458;
  wire[3:0] T22459;
  wire T22460;
  wire[46:0] twiddle4_1_493_imag;
  wire[46:0] T22461;
  wire[46:0] T22462;
  wire[46:0] T22463;
  wire[42:0] T22464;
  wire[42:0] T22465;
  wire[3:0] T22466;
  wire T22467;
  wire T22468;
  wire[46:0] T22469;
  wire[46:0] twiddle4_1_494_imag;
  wire[46:0] T22470;
  wire[46:0] T22471;
  wire[46:0] T22472;
  wire[42:0] T22473;
  wire[42:0] T22474;
  wire[3:0] T22475;
  wire T22476;
  wire[46:0] twiddle4_1_495_imag;
  wire[46:0] T22477;
  wire[46:0] T22478;
  wire[46:0] T22479;
  wire[42:0] T22480;
  wire[42:0] T22481;
  wire[3:0] T22482;
  wire T22483;
  wire T22484;
  wire T22485;
  wire T22486;
  wire T22487;
  wire[46:0] T22488;
  wire[46:0] T22489;
  wire[46:0] T22490;
  wire[46:0] T22491;
  wire[46:0] twiddle4_1_496_imag;
  wire[46:0] T22492;
  wire[46:0] T22493;
  wire[46:0] T22494;
  wire[42:0] T22495;
  wire[42:0] T22496;
  wire[3:0] T22497;
  wire T22498;
  wire[46:0] twiddle4_1_497_imag;
  wire[46:0] T22499;
  wire[46:0] T22500;
  wire[46:0] T22501;
  wire[42:0] T22502;
  wire[42:0] T22503;
  wire[3:0] T22504;
  wire T22505;
  wire T22506;
  wire[46:0] T22507;
  wire[46:0] twiddle4_1_498_imag;
  wire[46:0] T22508;
  wire[46:0] T22509;
  wire[46:0] T22510;
  wire[42:0] T22511;
  wire[42:0] T22512;
  wire[3:0] T22513;
  wire T22514;
  wire[46:0] twiddle4_1_499_imag;
  wire[46:0] T22515;
  wire[46:0] T22516;
  wire[46:0] T22517;
  wire[42:0] T22518;
  wire[42:0] T22519;
  wire[3:0] T22520;
  wire T22521;
  wire T22522;
  wire T22523;
  wire[46:0] T22524;
  wire[46:0] T22525;
  wire[46:0] twiddle4_1_500_imag;
  wire[46:0] T22526;
  wire[46:0] T22527;
  wire[46:0] T22528;
  wire[42:0] T22529;
  wire[42:0] T22530;
  wire[3:0] T22531;
  wire T22532;
  wire[46:0] twiddle4_1_501_imag;
  wire[46:0] T22533;
  wire[46:0] T22534;
  wire[46:0] T22535;
  wire[42:0] T22536;
  wire[42:0] T22537;
  wire[3:0] T22538;
  wire T22539;
  wire T22540;
  wire[46:0] T22541;
  wire[46:0] twiddle4_1_502_imag;
  wire[46:0] T22542;
  wire[46:0] T22543;
  wire[46:0] T22544;
  wire[41:0] T22545;
  wire[41:0] T22546;
  wire[4:0] T22547;
  wire T22548;
  wire[46:0] twiddle4_1_503_imag;
  wire[46:0] T22549;
  wire[46:0] T22550;
  wire[46:0] T22551;
  wire[41:0] T22552;
  wire[41:0] T22553;
  wire[4:0] T22554;
  wire T22555;
  wire T22556;
  wire T22557;
  wire T22558;
  wire[46:0] T22559;
  wire[46:0] T22560;
  wire[46:0] T22561;
  wire[46:0] twiddle4_1_504_imag;
  wire[46:0] T22562;
  wire[46:0] T22563;
  wire[46:0] T22564;
  wire[41:0] T22565;
  wire[41:0] T22566;
  wire[4:0] T22567;
  wire T22568;
  wire[46:0] twiddle4_1_505_imag;
  wire[46:0] T22569;
  wire[46:0] T22570;
  wire[46:0] T22571;
  wire[41:0] T22572;
  wire[41:0] T22573;
  wire[4:0] T22574;
  wire T22575;
  wire T22576;
  wire[46:0] T22577;
  wire[46:0] twiddle4_1_506_imag;
  wire[46:0] T22578;
  wire[46:0] T22579;
  wire[46:0] T22580;
  wire[41:0] T22581;
  wire[41:0] T22582;
  wire[4:0] T22583;
  wire T22584;
  wire[46:0] twiddle4_1_507_imag;
  wire[46:0] T22585;
  wire[46:0] T22586;
  wire[46:0] T22587;
  wire[40:0] T22588;
  wire[40:0] T22589;
  wire[5:0] T22590;
  wire T22591;
  wire T22592;
  wire T22593;
  wire[46:0] T22594;
  wire[46:0] T22595;
  wire[46:0] twiddle4_1_508_imag;
  wire[46:0] T22596;
  wire[46:0] T22597;
  wire[46:0] T22598;
  wire[40:0] T22599;
  wire[40:0] T22600;
  wire[5:0] T22601;
  wire T22602;
  wire[46:0] twiddle4_1_509_imag;
  wire[46:0] T22603;
  wire[46:0] T22604;
  wire[46:0] T22605;
  wire[40:0] T22606;
  wire[40:0] T22607;
  wire[5:0] T22608;
  wire T22609;
  wire T22610;
  wire[46:0] T22611;
  wire[46:0] twiddle4_1_510_imag;
  wire[46:0] T22612;
  wire[46:0] T22613;
  wire[46:0] T22614;
  wire[39:0] T22615;
  wire[39:0] T22616;
  wire[6:0] T22617;
  wire T22618;
  wire[46:0] twiddle4_1_511_imag;
  wire[46:0] T22619;
  wire[46:0] T22620;
  wire[46:0] T22621;
  wire[38:0] T22622;
  wire[38:0] T22623;
  wire[7:0] T22624;
  wire T22625;
  wire T22626;
  wire T22627;
  wire T22628;
  wire T22629;
  wire T22630;
  wire T22631;
  wire T22632;
  wire T22633;
  wire T22634;
  wire T22635;
  wire[15:0] T22636;
  wire[47:0] T22637;
  wire[47:0] T22638;
  wire[47:0] T22639;
  wire[47:0] T22640;
  wire[47:0] T22641;
  wire[47:0] T22642;
  wire[47:0] T22643;
  wire[47:0] T22644;
  wire[47:0] T22645;
  wire[47:0] twiddle4_1_0_real;
  wire[47:0] T22646;
  wire[16:0] T22647;
  wire[16:0] T22648;
  wire[30:0] T22649;
  wire T22650;
  wire[47:0] T22651;
  wire[47:0] T22652;
  wire[47:0] T22653;
  wire[46:0] twiddle4_1_1_real;
  wire[46:0] T22654;
  wire[38:0] T22655;
  wire[38:0] T22656;
  wire[7:0] T22657;
  wire T22658;
  wire[46:0] T22659;
  wire[46:0] T22660;
  wire T22661;
  wire T22662;
  wire[47:0] T22663;
  wire[46:0] T22664;
  wire[46:0] twiddle4_1_2_real;
  wire[46:0] T22665;
  wire[39:0] T22666;
  wire[39:0] T22667;
  wire[6:0] T22668;
  wire T22669;
  wire[46:0] T22670;
  wire[46:0] T22671;
  wire[46:0] twiddle4_1_3_real;
  wire[46:0] T22672;
  wire[40:0] T22673;
  wire[40:0] T22674;
  wire[5:0] T22675;
  wire T22676;
  wire[46:0] T22677;
  wire[46:0] T22678;
  wire T22679;
  wire T22680;
  wire T22681;
  wire[47:0] T22682;
  wire[46:0] T22683;
  wire[46:0] T22684;
  wire[46:0] twiddle4_1_4_real;
  wire[46:0] T22685;
  wire[40:0] T22686;
  wire[40:0] T22687;
  wire[5:0] T22688;
  wire T22689;
  wire[46:0] T22690;
  wire[46:0] T22691;
  wire[46:0] twiddle4_1_5_real;
  wire[46:0] T22692;
  wire[40:0] T22693;
  wire[40:0] T22694;
  wire[5:0] T22695;
  wire T22696;
  wire[46:0] T22697;
  wire[46:0] T22698;
  wire T22699;
  wire[46:0] T22700;
  wire[46:0] twiddle4_1_6_real;
  wire[46:0] T22701;
  wire[41:0] T22702;
  wire[41:0] T22703;
  wire[4:0] T22704;
  wire T22705;
  wire[46:0] T22706;
  wire[46:0] T22707;
  wire[46:0] twiddle4_1_7_real;
  wire[46:0] T22708;
  wire[41:0] T22709;
  wire[41:0] T22710;
  wire[4:0] T22711;
  wire T22712;
  wire[46:0] T22713;
  wire[46:0] T22714;
  wire T22715;
  wire T22716;
  wire T22717;
  wire T22718;
  wire[47:0] T22719;
  wire[46:0] T22720;
  wire[46:0] T22721;
  wire[46:0] T22722;
  wire[46:0] twiddle4_1_8_real;
  wire[46:0] T22723;
  wire[41:0] T22724;
  wire[41:0] T22725;
  wire[4:0] T22726;
  wire T22727;
  wire[46:0] T22728;
  wire[46:0] T22729;
  wire[46:0] twiddle4_1_9_real;
  wire[46:0] T22730;
  wire[41:0] T22731;
  wire[41:0] T22732;
  wire[4:0] T22733;
  wire T22734;
  wire[46:0] T22735;
  wire[46:0] T22736;
  wire T22737;
  wire[46:0] T22738;
  wire[46:0] twiddle4_1_10_real;
  wire[46:0] T22739;
  wire[41:0] T22740;
  wire[41:0] T22741;
  wire[4:0] T22742;
  wire T22743;
  wire[46:0] T22744;
  wire[46:0] T22745;
  wire[46:0] twiddle4_1_11_real;
  wire[46:0] T22746;
  wire[42:0] T22747;
  wire[42:0] T22748;
  wire[3:0] T22749;
  wire T22750;
  wire[46:0] T22751;
  wire[46:0] T22752;
  wire T22753;
  wire T22754;
  wire[46:0] T22755;
  wire[46:0] T22756;
  wire[46:0] twiddle4_1_12_real;
  wire[46:0] T22757;
  wire[42:0] T22758;
  wire[42:0] T22759;
  wire[3:0] T22760;
  wire T22761;
  wire[46:0] T22762;
  wire[46:0] T22763;
  wire[46:0] twiddle4_1_13_real;
  wire[46:0] T22764;
  wire[42:0] T22765;
  wire[42:0] T22766;
  wire[3:0] T22767;
  wire T22768;
  wire[46:0] T22769;
  wire[46:0] T22770;
  wire T22771;
  wire[46:0] T22772;
  wire[46:0] twiddle4_1_14_real;
  wire[46:0] T22773;
  wire[42:0] T22774;
  wire[42:0] T22775;
  wire[3:0] T22776;
  wire T22777;
  wire[46:0] T22778;
  wire[46:0] T22779;
  wire[46:0] twiddle4_1_15_real;
  wire[46:0] T22780;
  wire[42:0] T22781;
  wire[42:0] T22782;
  wire[3:0] T22783;
  wire T22784;
  wire[46:0] T22785;
  wire[46:0] T22786;
  wire T22787;
  wire T22788;
  wire T22789;
  wire T22790;
  wire T22791;
  wire[47:0] T22792;
  wire[46:0] T22793;
  wire[46:0] T22794;
  wire[46:0] T22795;
  wire[46:0] T22796;
  wire[46:0] twiddle4_1_16_real;
  wire[46:0] T22797;
  wire[42:0] T22798;
  wire[42:0] T22799;
  wire[3:0] T22800;
  wire T22801;
  wire[46:0] T22802;
  wire[46:0] T22803;
  wire[46:0] twiddle4_1_17_real;
  wire[46:0] T22804;
  wire[42:0] T22805;
  wire[42:0] T22806;
  wire[3:0] T22807;
  wire T22808;
  wire[46:0] T22809;
  wire[46:0] T22810;
  wire T22811;
  wire[46:0] T22812;
  wire[46:0] twiddle4_1_18_real;
  wire[46:0] T22813;
  wire[42:0] T22814;
  wire[42:0] T22815;
  wire[3:0] T22816;
  wire T22817;
  wire[46:0] T22818;
  wire[46:0] T22819;
  wire[46:0] twiddle4_1_19_real;
  wire[46:0] T22820;
  wire[42:0] T22821;
  wire[42:0] T22822;
  wire[3:0] T22823;
  wire T22824;
  wire[46:0] T22825;
  wire[46:0] T22826;
  wire T22827;
  wire T22828;
  wire[46:0] T22829;
  wire[46:0] T22830;
  wire[46:0] twiddle4_1_20_real;
  wire[46:0] T22831;
  wire[42:0] T22832;
  wire[42:0] T22833;
  wire[3:0] T22834;
  wire T22835;
  wire[46:0] T22836;
  wire[46:0] T22837;
  wire[46:0] twiddle4_1_21_real;
  wire[46:0] T22838;
  wire[43:0] T22839;
  wire[43:0] T22840;
  wire[2:0] T22841;
  wire T22842;
  wire[46:0] T22843;
  wire[46:0] T22844;
  wire T22845;
  wire[46:0] T22846;
  wire[46:0] twiddle4_1_22_real;
  wire[46:0] T22847;
  wire[43:0] T22848;
  wire[43:0] T22849;
  wire[2:0] T22850;
  wire T22851;
  wire[46:0] T22852;
  wire[46:0] T22853;
  wire[46:0] twiddle4_1_23_real;
  wire[46:0] T22854;
  wire[43:0] T22855;
  wire[43:0] T22856;
  wire[2:0] T22857;
  wire T22858;
  wire[46:0] T22859;
  wire[46:0] T22860;
  wire T22861;
  wire T22862;
  wire T22863;
  wire[46:0] T22864;
  wire[46:0] T22865;
  wire[46:0] T22866;
  wire[46:0] twiddle4_1_24_real;
  wire[46:0] T22867;
  wire[43:0] T22868;
  wire[43:0] T22869;
  wire[2:0] T22870;
  wire T22871;
  wire[46:0] T22872;
  wire[46:0] T22873;
  wire[46:0] twiddle4_1_25_real;
  wire[46:0] T22874;
  wire[43:0] T22875;
  wire[43:0] T22876;
  wire[2:0] T22877;
  wire T22878;
  wire[46:0] T22879;
  wire[46:0] T22880;
  wire T22881;
  wire[46:0] T22882;
  wire[46:0] twiddle4_1_26_real;
  wire[46:0] T22883;
  wire[43:0] T22884;
  wire[43:0] T22885;
  wire[2:0] T22886;
  wire T22887;
  wire[46:0] T22888;
  wire[46:0] T22889;
  wire[46:0] twiddle4_1_27_real;
  wire[46:0] T22890;
  wire[43:0] T22891;
  wire[43:0] T22892;
  wire[2:0] T22893;
  wire T22894;
  wire[46:0] T22895;
  wire[46:0] T22896;
  wire T22897;
  wire T22898;
  wire[46:0] T22899;
  wire[46:0] T22900;
  wire[46:0] twiddle4_1_28_real;
  wire[46:0] T22901;
  wire[43:0] T22902;
  wire[43:0] T22903;
  wire[2:0] T22904;
  wire T22905;
  wire[46:0] T22906;
  wire[46:0] T22907;
  wire[46:0] twiddle4_1_29_real;
  wire[46:0] T22908;
  wire[43:0] T22909;
  wire[43:0] T22910;
  wire[2:0] T22911;
  wire T22912;
  wire[46:0] T22913;
  wire[46:0] T22914;
  wire T22915;
  wire[46:0] T22916;
  wire[46:0] twiddle4_1_30_real;
  wire[46:0] T22917;
  wire[43:0] T22918;
  wire[43:0] T22919;
  wire[2:0] T22920;
  wire T22921;
  wire[46:0] T22922;
  wire[46:0] T22923;
  wire[46:0] twiddle4_1_31_real;
  wire[46:0] T22924;
  wire[43:0] T22925;
  wire[43:0] T22926;
  wire[2:0] T22927;
  wire T22928;
  wire[46:0] T22929;
  wire[46:0] T22930;
  wire T22931;
  wire T22932;
  wire T22933;
  wire T22934;
  wire T22935;
  wire T22936;
  wire[47:0] T22937;
  wire[46:0] T22938;
  wire[46:0] T22939;
  wire[46:0] T22940;
  wire[46:0] T22941;
  wire[46:0] T22942;
  wire[46:0] twiddle4_1_32_real;
  wire[46:0] T22943;
  wire[43:0] T22944;
  wire[43:0] T22945;
  wire[2:0] T22946;
  wire T22947;
  wire[46:0] T22948;
  wire[46:0] T22949;
  wire[46:0] twiddle4_1_33_real;
  wire[46:0] T22950;
  wire[43:0] T22951;
  wire[43:0] T22952;
  wire[2:0] T22953;
  wire T22954;
  wire[46:0] T22955;
  wire[46:0] T22956;
  wire T22957;
  wire[46:0] T22958;
  wire[46:0] twiddle4_1_34_real;
  wire[46:0] T22959;
  wire[43:0] T22960;
  wire[43:0] T22961;
  wire[2:0] T22962;
  wire T22963;
  wire[46:0] T22964;
  wire[46:0] T22965;
  wire[46:0] twiddle4_1_35_real;
  wire[46:0] T22966;
  wire[43:0] T22967;
  wire[43:0] T22968;
  wire[2:0] T22969;
  wire T22970;
  wire[46:0] T22971;
  wire[46:0] T22972;
  wire T22973;
  wire T22974;
  wire[46:0] T22975;
  wire[46:0] T22976;
  wire[46:0] twiddle4_1_36_real;
  wire[46:0] T22977;
  wire[43:0] T22978;
  wire[43:0] T22979;
  wire[2:0] T22980;
  wire T22981;
  wire[46:0] T22982;
  wire[46:0] T22983;
  wire[46:0] twiddle4_1_37_real;
  wire[46:0] T22984;
  wire[43:0] T22985;
  wire[43:0] T22986;
  wire[2:0] T22987;
  wire T22988;
  wire[46:0] T22989;
  wire[46:0] T22990;
  wire T22991;
  wire[46:0] T22992;
  wire[46:0] twiddle4_1_38_real;
  wire[46:0] T22993;
  wire[43:0] T22994;
  wire[43:0] T22995;
  wire[2:0] T22996;
  wire T22997;
  wire[46:0] T22998;
  wire[46:0] T22999;
  wire[46:0] twiddle4_1_39_real;
  wire[46:0] T23000;
  wire[43:0] T23001;
  wire[43:0] T23002;
  wire[2:0] T23003;
  wire T23004;
  wire[46:0] T23005;
  wire[46:0] T23006;
  wire T23007;
  wire T23008;
  wire T23009;
  wire[46:0] T23010;
  wire[46:0] T23011;
  wire[46:0] T23012;
  wire[46:0] twiddle4_1_40_real;
  wire[46:0] T23013;
  wire[43:0] T23014;
  wire[43:0] T23015;
  wire[2:0] T23016;
  wire T23017;
  wire[46:0] T23018;
  wire[46:0] T23019;
  wire[46:0] twiddle4_1_41_real;
  wire[46:0] T23020;
  wire[44:0] T23021;
  wire[44:0] T23022;
  wire[1:0] T23023;
  wire T23024;
  wire[46:0] T23025;
  wire[46:0] T23026;
  wire T23027;
  wire[46:0] T23028;
  wire[46:0] twiddle4_1_42_real;
  wire[46:0] T23029;
  wire[44:0] T23030;
  wire[44:0] T23031;
  wire[1:0] T23032;
  wire T23033;
  wire[46:0] T23034;
  wire[46:0] T23035;
  wire[46:0] twiddle4_1_43_real;
  wire[46:0] T23036;
  wire[44:0] T23037;
  wire[44:0] T23038;
  wire[1:0] T23039;
  wire T23040;
  wire[46:0] T23041;
  wire[46:0] T23042;
  wire T23043;
  wire T23044;
  wire[46:0] T23045;
  wire[46:0] T23046;
  wire[46:0] twiddle4_1_44_real;
  wire[46:0] T23047;
  wire[44:0] T23048;
  wire[44:0] T23049;
  wire[1:0] T23050;
  wire T23051;
  wire[46:0] T23052;
  wire[46:0] T23053;
  wire[46:0] twiddle4_1_45_real;
  wire[46:0] T23054;
  wire[44:0] T23055;
  wire[44:0] T23056;
  wire[1:0] T23057;
  wire T23058;
  wire[46:0] T23059;
  wire[46:0] T23060;
  wire T23061;
  wire[46:0] T23062;
  wire[46:0] twiddle4_1_46_real;
  wire[46:0] T23063;
  wire[44:0] T23064;
  wire[44:0] T23065;
  wire[1:0] T23066;
  wire T23067;
  wire[46:0] T23068;
  wire[46:0] T23069;
  wire[46:0] twiddle4_1_47_real;
  wire[46:0] T23070;
  wire[44:0] T23071;
  wire[44:0] T23072;
  wire[1:0] T23073;
  wire T23074;
  wire[46:0] T23075;
  wire[46:0] T23076;
  wire T23077;
  wire T23078;
  wire T23079;
  wire T23080;
  wire[46:0] T23081;
  wire[46:0] T23082;
  wire[46:0] T23083;
  wire[46:0] T23084;
  wire[46:0] twiddle4_1_48_real;
  wire[46:0] T23085;
  wire[44:0] T23086;
  wire[44:0] T23087;
  wire[1:0] T23088;
  wire T23089;
  wire[46:0] T23090;
  wire[46:0] T23091;
  wire[46:0] twiddle4_1_49_real;
  wire[46:0] T23092;
  wire[44:0] T23093;
  wire[44:0] T23094;
  wire[1:0] T23095;
  wire T23096;
  wire[46:0] T23097;
  wire[46:0] T23098;
  wire T23099;
  wire[46:0] T23100;
  wire[46:0] twiddle4_1_50_real;
  wire[46:0] T23101;
  wire[44:0] T23102;
  wire[44:0] T23103;
  wire[1:0] T23104;
  wire T23105;
  wire[46:0] T23106;
  wire[46:0] T23107;
  wire[46:0] twiddle4_1_51_real;
  wire[46:0] T23108;
  wire[44:0] T23109;
  wire[44:0] T23110;
  wire[1:0] T23111;
  wire T23112;
  wire[46:0] T23113;
  wire[46:0] T23114;
  wire T23115;
  wire T23116;
  wire[46:0] T23117;
  wire[46:0] T23118;
  wire[46:0] twiddle4_1_52_real;
  wire[46:0] T23119;
  wire[44:0] T23120;
  wire[44:0] T23121;
  wire[1:0] T23122;
  wire T23123;
  wire[46:0] T23124;
  wire[46:0] T23125;
  wire[46:0] twiddle4_1_53_real;
  wire[46:0] T23126;
  wire[44:0] T23127;
  wire[44:0] T23128;
  wire[1:0] T23129;
  wire T23130;
  wire[46:0] T23131;
  wire[46:0] T23132;
  wire T23133;
  wire[46:0] T23134;
  wire[46:0] twiddle4_1_54_real;
  wire[46:0] T23135;
  wire[44:0] T23136;
  wire[44:0] T23137;
  wire[1:0] T23138;
  wire T23139;
  wire[46:0] T23140;
  wire[46:0] T23141;
  wire[46:0] twiddle4_1_55_real;
  wire[46:0] T23142;
  wire[44:0] T23143;
  wire[44:0] T23144;
  wire[1:0] T23145;
  wire T23146;
  wire[46:0] T23147;
  wire[46:0] T23148;
  wire T23149;
  wire T23150;
  wire T23151;
  wire[46:0] T23152;
  wire[46:0] T23153;
  wire[46:0] T23154;
  wire[46:0] twiddle4_1_56_real;
  wire[46:0] T23155;
  wire[44:0] T23156;
  wire[44:0] T23157;
  wire[1:0] T23158;
  wire T23159;
  wire[46:0] T23160;
  wire[46:0] T23161;
  wire[46:0] twiddle4_1_57_real;
  wire[46:0] T23162;
  wire[44:0] T23163;
  wire[44:0] T23164;
  wire[1:0] T23165;
  wire T23166;
  wire[46:0] T23167;
  wire[46:0] T23168;
  wire T23169;
  wire[46:0] T23170;
  wire[46:0] twiddle4_1_58_real;
  wire[46:0] T23171;
  wire[44:0] T23172;
  wire[44:0] T23173;
  wire[1:0] T23174;
  wire T23175;
  wire[46:0] T23176;
  wire[46:0] T23177;
  wire[46:0] twiddle4_1_59_real;
  wire[46:0] T23178;
  wire[44:0] T23179;
  wire[44:0] T23180;
  wire[1:0] T23181;
  wire T23182;
  wire[46:0] T23183;
  wire[46:0] T23184;
  wire T23185;
  wire T23186;
  wire[46:0] T23187;
  wire[46:0] T23188;
  wire[46:0] twiddle4_1_60_real;
  wire[46:0] T23189;
  wire[44:0] T23190;
  wire[44:0] T23191;
  wire[1:0] T23192;
  wire T23193;
  wire[46:0] T23194;
  wire[46:0] T23195;
  wire[46:0] twiddle4_1_61_real;
  wire[46:0] T23196;
  wire[44:0] T23197;
  wire[44:0] T23198;
  wire[1:0] T23199;
  wire T23200;
  wire[46:0] T23201;
  wire[46:0] T23202;
  wire T23203;
  wire[46:0] T23204;
  wire[46:0] twiddle4_1_62_real;
  wire[46:0] T23205;
  wire[44:0] T23206;
  wire[44:0] T23207;
  wire[1:0] T23208;
  wire T23209;
  wire[46:0] T23210;
  wire[46:0] T23211;
  wire[46:0] twiddle4_1_63_real;
  wire[46:0] T23212;
  wire[44:0] T23213;
  wire[44:0] T23214;
  wire[1:0] T23215;
  wire T23216;
  wire[46:0] T23217;
  wire[46:0] T23218;
  wire T23219;
  wire T23220;
  wire T23221;
  wire T23222;
  wire T23223;
  wire T23224;
  wire T23225;
  wire[47:0] T23226;
  wire[46:0] T23227;
  wire[46:0] T23228;
  wire[46:0] T23229;
  wire[46:0] T23230;
  wire[46:0] T23231;
  wire[46:0] T23232;
  wire[46:0] twiddle4_1_64_real;
  wire[46:0] T23233;
  wire[44:0] T23234;
  wire[44:0] T23235;
  wire[1:0] T23236;
  wire T23237;
  wire[46:0] T23238;
  wire[46:0] T23239;
  wire[46:0] twiddle4_1_65_real;
  wire[46:0] T23240;
  wire[44:0] T23241;
  wire[44:0] T23242;
  wire[1:0] T23243;
  wire T23244;
  wire[46:0] T23245;
  wire[46:0] T23246;
  wire T23247;
  wire[46:0] T23248;
  wire[46:0] twiddle4_1_66_real;
  wire[46:0] T23249;
  wire[44:0] T23250;
  wire[44:0] T23251;
  wire[1:0] T23252;
  wire T23253;
  wire[46:0] T23254;
  wire[46:0] T23255;
  wire[46:0] twiddle4_1_67_real;
  wire[46:0] T23256;
  wire[44:0] T23257;
  wire[44:0] T23258;
  wire[1:0] T23259;
  wire T23260;
  wire[46:0] T23261;
  wire[46:0] T23262;
  wire T23263;
  wire T23264;
  wire[46:0] T23265;
  wire[46:0] T23266;
  wire[46:0] twiddle4_1_68_real;
  wire[46:0] T23267;
  wire[44:0] T23268;
  wire[44:0] T23269;
  wire[1:0] T23270;
  wire T23271;
  wire[46:0] T23272;
  wire[46:0] T23273;
  wire[46:0] twiddle4_1_69_real;
  wire[46:0] T23274;
  wire[44:0] T23275;
  wire[44:0] T23276;
  wire[1:0] T23277;
  wire T23278;
  wire[46:0] T23279;
  wire[46:0] T23280;
  wire T23281;
  wire[46:0] T23282;
  wire[46:0] twiddle4_1_70_real;
  wire[46:0] T23283;
  wire[44:0] T23284;
  wire[44:0] T23285;
  wire[1:0] T23286;
  wire T23287;
  wire[46:0] T23288;
  wire[46:0] T23289;
  wire[46:0] twiddle4_1_71_real;
  wire[46:0] T23290;
  wire[44:0] T23291;
  wire[44:0] T23292;
  wire[1:0] T23293;
  wire T23294;
  wire[46:0] T23295;
  wire[46:0] T23296;
  wire T23297;
  wire T23298;
  wire T23299;
  wire[46:0] T23300;
  wire[46:0] T23301;
  wire[46:0] T23302;
  wire[46:0] twiddle4_1_72_real;
  wire[46:0] T23303;
  wire[44:0] T23304;
  wire[44:0] T23305;
  wire[1:0] T23306;
  wire T23307;
  wire[46:0] T23308;
  wire[46:0] T23309;
  wire[46:0] twiddle4_1_73_real;
  wire[46:0] T23310;
  wire[44:0] T23311;
  wire[44:0] T23312;
  wire[1:0] T23313;
  wire T23314;
  wire[46:0] T23315;
  wire[46:0] T23316;
  wire T23317;
  wire[46:0] T23318;
  wire[46:0] twiddle4_1_74_real;
  wire[46:0] T23319;
  wire[44:0] T23320;
  wire[44:0] T23321;
  wire[1:0] T23322;
  wire T23323;
  wire[46:0] T23324;
  wire[46:0] T23325;
  wire[46:0] twiddle4_1_75_real;
  wire[46:0] T23326;
  wire[44:0] T23327;
  wire[44:0] T23328;
  wire[1:0] T23329;
  wire T23330;
  wire[46:0] T23331;
  wire[46:0] T23332;
  wire T23333;
  wire T23334;
  wire[46:0] T23335;
  wire[46:0] T23336;
  wire[46:0] twiddle4_1_76_real;
  wire[46:0] T23337;
  wire[44:0] T23338;
  wire[44:0] T23339;
  wire[1:0] T23340;
  wire T23341;
  wire[46:0] T23342;
  wire[46:0] T23343;
  wire[46:0] twiddle4_1_77_real;
  wire[46:0] T23344;
  wire[44:0] T23345;
  wire[44:0] T23346;
  wire[1:0] T23347;
  wire T23348;
  wire[46:0] T23349;
  wire[46:0] T23350;
  wire T23351;
  wire[46:0] T23352;
  wire[46:0] twiddle4_1_78_real;
  wire[46:0] T23353;
  wire[44:0] T23354;
  wire[44:0] T23355;
  wire[1:0] T23356;
  wire T23357;
  wire[46:0] T23358;
  wire[46:0] T23359;
  wire[46:0] twiddle4_1_79_real;
  wire[46:0] T23360;
  wire[44:0] T23361;
  wire[44:0] T23362;
  wire[1:0] T23363;
  wire T23364;
  wire[46:0] T23365;
  wire[46:0] T23366;
  wire T23367;
  wire T23368;
  wire T23369;
  wire T23370;
  wire[46:0] T23371;
  wire[46:0] T23372;
  wire[46:0] T23373;
  wire[46:0] T23374;
  wire[46:0] twiddle4_1_80_real;
  wire[46:0] T23375;
  wire[44:0] T23376;
  wire[44:0] T23377;
  wire[1:0] T23378;
  wire T23379;
  wire[46:0] T23380;
  wire[46:0] T23381;
  wire[46:0] twiddle4_1_81_real;
  wire[46:0] T23382;
  wire[44:0] T23383;
  wire[44:0] T23384;
  wire[1:0] T23385;
  wire T23386;
  wire[46:0] T23387;
  wire[46:0] T23388;
  wire T23389;
  wire[46:0] T23390;
  wire[46:0] twiddle4_1_82_real;
  wire[46:0] T23391;
  wire[44:0] T23392;
  wire[44:0] T23393;
  wire[1:0] T23394;
  wire T23395;
  wire[46:0] T23396;
  wire[46:0] T23397;
  wire[46:0] twiddle4_1_83_real;
  wire[46:0] T23398;
  wire[45:0] T23399;
  wire[45:0] T23400;
  wire T23401;
  wire[46:0] T23402;
  wire[46:0] T23403;
  wire T23404;
  wire T23405;
  wire[46:0] T23406;
  wire[46:0] T23407;
  wire[46:0] twiddle4_1_84_real;
  wire[46:0] T23408;
  wire[45:0] T23409;
  wire[45:0] T23410;
  wire T23411;
  wire[46:0] T23412;
  wire[46:0] T23413;
  wire[46:0] twiddle4_1_85_real;
  wire[46:0] T23414;
  wire[45:0] T23415;
  wire[45:0] T23416;
  wire T23417;
  wire[46:0] T23418;
  wire[46:0] T23419;
  wire T23420;
  wire[46:0] T23421;
  wire[46:0] twiddle4_1_86_real;
  wire[46:0] T23422;
  wire[45:0] T23423;
  wire[45:0] T23424;
  wire T23425;
  wire[46:0] T23426;
  wire[46:0] T23427;
  wire[46:0] twiddle4_1_87_real;
  wire[46:0] T23428;
  wire[45:0] T23429;
  wire[45:0] T23430;
  wire T23431;
  wire[46:0] T23432;
  wire[46:0] T23433;
  wire T23434;
  wire T23435;
  wire T23436;
  wire[46:0] T23437;
  wire[46:0] T23438;
  wire[46:0] T23439;
  wire[46:0] twiddle4_1_88_real;
  wire[46:0] T23440;
  wire[45:0] T23441;
  wire[45:0] T23442;
  wire T23443;
  wire[46:0] T23444;
  wire[46:0] T23445;
  wire[46:0] twiddle4_1_89_real;
  wire[46:0] T23446;
  wire[45:0] T23447;
  wire[45:0] T23448;
  wire T23449;
  wire[46:0] T23450;
  wire[46:0] T23451;
  wire T23452;
  wire[46:0] T23453;
  wire[46:0] twiddle4_1_90_real;
  wire[46:0] T23454;
  wire[45:0] T23455;
  wire[45:0] T23456;
  wire T23457;
  wire[46:0] T23458;
  wire[46:0] T23459;
  wire[46:0] twiddle4_1_91_real;
  wire[46:0] T23460;
  wire[45:0] T23461;
  wire[45:0] T23462;
  wire T23463;
  wire[46:0] T23464;
  wire[46:0] T23465;
  wire T23466;
  wire T23467;
  wire[46:0] T23468;
  wire[46:0] T23469;
  wire[46:0] twiddle4_1_92_real;
  wire[46:0] T23470;
  wire[45:0] T23471;
  wire[45:0] T23472;
  wire T23473;
  wire[46:0] T23474;
  wire[46:0] T23475;
  wire[46:0] twiddle4_1_93_real;
  wire[46:0] T23476;
  wire[45:0] T23477;
  wire[45:0] T23478;
  wire T23479;
  wire[46:0] T23480;
  wire[46:0] T23481;
  wire T23482;
  wire[46:0] T23483;
  wire[46:0] twiddle4_1_94_real;
  wire[46:0] T23484;
  wire[45:0] T23485;
  wire[45:0] T23486;
  wire T23487;
  wire[46:0] T23488;
  wire[46:0] T23489;
  wire[46:0] twiddle4_1_95_real;
  wire[46:0] T23490;
  wire[45:0] T23491;
  wire[45:0] T23492;
  wire T23493;
  wire[46:0] T23494;
  wire[46:0] T23495;
  wire T23496;
  wire T23497;
  wire T23498;
  wire T23499;
  wire T23500;
  wire[46:0] T23501;
  wire[46:0] T23502;
  wire[46:0] T23503;
  wire[46:0] T23504;
  wire[46:0] T23505;
  wire[46:0] twiddle4_1_96_real;
  wire[46:0] T23506;
  wire[45:0] T23507;
  wire[45:0] T23508;
  wire T23509;
  wire[46:0] T23510;
  wire[46:0] T23511;
  wire[46:0] twiddle4_1_97_real;
  wire[46:0] T23512;
  wire[45:0] T23513;
  wire[45:0] T23514;
  wire T23515;
  wire[46:0] T23516;
  wire[46:0] T23517;
  wire T23518;
  wire[46:0] T23519;
  wire[46:0] twiddle4_1_98_real;
  wire[46:0] T23520;
  wire[45:0] T23521;
  wire[45:0] T23522;
  wire T23523;
  wire[46:0] T23524;
  wire[46:0] T23525;
  wire[46:0] twiddle4_1_99_real;
  wire[46:0] T23526;
  wire[45:0] T23527;
  wire[45:0] T23528;
  wire T23529;
  wire[46:0] T23530;
  wire[46:0] T23531;
  wire T23532;
  wire T23533;
  wire[46:0] T23534;
  wire[46:0] T23535;
  wire[46:0] twiddle4_1_100_real;
  wire[46:0] T23536;
  wire[45:0] T23537;
  wire[45:0] T23538;
  wire T23539;
  wire[46:0] T23540;
  wire[46:0] T23541;
  wire[46:0] twiddle4_1_101_real;
  wire[46:0] T23542;
  wire[45:0] T23543;
  wire[45:0] T23544;
  wire T23545;
  wire[46:0] T23546;
  wire[46:0] T23547;
  wire T23548;
  wire[46:0] T23549;
  wire[46:0] twiddle4_1_102_real;
  wire[46:0] T23550;
  wire[45:0] T23551;
  wire[45:0] T23552;
  wire T23553;
  wire[46:0] T23554;
  wire[46:0] T23555;
  wire[46:0] twiddle4_1_103_real;
  wire[46:0] T23556;
  wire[45:0] T23557;
  wire[45:0] T23558;
  wire T23559;
  wire[46:0] T23560;
  wire[46:0] T23561;
  wire T23562;
  wire T23563;
  wire T23564;
  wire[46:0] T23565;
  wire[46:0] T23566;
  wire[46:0] T23567;
  wire[46:0] twiddle4_1_104_real;
  wire[46:0] T23568;
  wire[45:0] T23569;
  wire[45:0] T23570;
  wire T23571;
  wire[46:0] T23572;
  wire[46:0] T23573;
  wire[46:0] twiddle4_1_105_real;
  wire[46:0] T23574;
  wire[45:0] T23575;
  wire[45:0] T23576;
  wire T23577;
  wire[46:0] T23578;
  wire[46:0] T23579;
  wire T23580;
  wire[46:0] T23581;
  wire[46:0] twiddle4_1_106_real;
  wire[46:0] T23582;
  wire[45:0] T23583;
  wire[45:0] T23584;
  wire T23585;
  wire[46:0] T23586;
  wire[46:0] T23587;
  wire[46:0] twiddle4_1_107_real;
  wire[46:0] T23588;
  wire[45:0] T23589;
  wire[45:0] T23590;
  wire T23591;
  wire[46:0] T23592;
  wire[46:0] T23593;
  wire T23594;
  wire T23595;
  wire[46:0] T23596;
  wire[46:0] T23597;
  wire[46:0] twiddle4_1_108_real;
  wire[46:0] T23598;
  wire[45:0] T23599;
  wire[45:0] T23600;
  wire T23601;
  wire[46:0] T23602;
  wire[46:0] T23603;
  wire[46:0] twiddle4_1_109_real;
  wire[46:0] T23604;
  wire[45:0] T23605;
  wire[45:0] T23606;
  wire T23607;
  wire[46:0] T23608;
  wire[46:0] T23609;
  wire T23610;
  wire[46:0] T23611;
  wire[46:0] twiddle4_1_110_real;
  wire[46:0] T23612;
  wire[45:0] T23613;
  wire[45:0] T23614;
  wire T23615;
  wire[46:0] T23616;
  wire[46:0] T23617;
  wire[46:0] twiddle4_1_111_real;
  wire[46:0] T23618;
  wire[45:0] T23619;
  wire[45:0] T23620;
  wire T23621;
  wire[46:0] T23622;
  wire[46:0] T23623;
  wire T23624;
  wire T23625;
  wire T23626;
  wire T23627;
  wire[46:0] T23628;
  wire[46:0] T23629;
  wire[46:0] T23630;
  wire[46:0] T23631;
  wire[46:0] twiddle4_1_112_real;
  wire[46:0] T23632;
  wire[45:0] T23633;
  wire[45:0] T23634;
  wire T23635;
  wire[46:0] T23636;
  wire[46:0] T23637;
  wire[46:0] twiddle4_1_113_real;
  wire[46:0] T23638;
  wire[45:0] T23639;
  wire[45:0] T23640;
  wire T23641;
  wire[46:0] T23642;
  wire[46:0] T23643;
  wire T23644;
  wire[46:0] T23645;
  wire[46:0] twiddle4_1_114_real;
  wire[46:0] T23646;
  wire[45:0] T23647;
  wire[45:0] T23648;
  wire T23649;
  wire[46:0] T23650;
  wire[46:0] T23651;
  wire[46:0] twiddle4_1_115_real;
  wire[46:0] T23652;
  wire[45:0] T23653;
  wire[45:0] T23654;
  wire T23655;
  wire[46:0] T23656;
  wire[46:0] T23657;
  wire T23658;
  wire T23659;
  wire[46:0] T23660;
  wire[46:0] T23661;
  wire[46:0] twiddle4_1_116_real;
  wire[46:0] T23662;
  wire[45:0] T23663;
  wire[45:0] T23664;
  wire T23665;
  wire[46:0] T23666;
  wire[46:0] T23667;
  wire[46:0] twiddle4_1_117_real;
  wire[46:0] T23668;
  wire[45:0] T23669;
  wire[45:0] T23670;
  wire T23671;
  wire[46:0] T23672;
  wire[46:0] T23673;
  wire T23674;
  wire[46:0] T23675;
  wire[46:0] twiddle4_1_118_real;
  wire[46:0] T23676;
  wire[45:0] T23677;
  wire[45:0] T23678;
  wire T23679;
  wire[46:0] T23680;
  wire[46:0] T23681;
  wire[46:0] twiddle4_1_119_real;
  wire[46:0] T23682;
  wire[45:0] T23683;
  wire[45:0] T23684;
  wire T23685;
  wire[46:0] T23686;
  wire[46:0] T23687;
  wire T23688;
  wire T23689;
  wire T23690;
  wire[46:0] T23691;
  wire[46:0] T23692;
  wire[46:0] T23693;
  wire[46:0] twiddle4_1_120_real;
  wire[46:0] T23694;
  wire[45:0] T23695;
  wire[45:0] T23696;
  wire T23697;
  wire[46:0] T23698;
  wire[46:0] T23699;
  wire[46:0] twiddle4_1_121_real;
  wire[46:0] T23700;
  wire[45:0] T23701;
  wire[45:0] T23702;
  wire T23703;
  wire[46:0] T23704;
  wire[46:0] T23705;
  wire T23706;
  wire[46:0] T23707;
  wire[46:0] twiddle4_1_122_real;
  wire[46:0] T23708;
  wire[45:0] T23709;
  wire[45:0] T23710;
  wire T23711;
  wire[46:0] T23712;
  wire[46:0] T23713;
  wire[46:0] twiddle4_1_123_real;
  wire[46:0] T23714;
  wire[45:0] T23715;
  wire[45:0] T23716;
  wire T23717;
  wire[46:0] T23718;
  wire[46:0] T23719;
  wire T23720;
  wire T23721;
  wire[46:0] T23722;
  wire[46:0] T23723;
  wire[46:0] twiddle4_1_124_real;
  wire[46:0] T23724;
  wire[45:0] T23725;
  wire[45:0] T23726;
  wire T23727;
  wire[46:0] T23728;
  wire[46:0] T23729;
  wire[46:0] twiddle4_1_125_real;
  wire[46:0] T23730;
  wire[45:0] T23731;
  wire[45:0] T23732;
  wire T23733;
  wire[46:0] T23734;
  wire[46:0] T23735;
  wire T23736;
  wire[46:0] T23737;
  wire[46:0] twiddle4_1_126_real;
  wire[46:0] T23738;
  wire[45:0] T23739;
  wire[45:0] T23740;
  wire T23741;
  wire[46:0] T23742;
  wire[46:0] T23743;
  wire[46:0] twiddle4_1_127_real;
  wire[46:0] T23744;
  wire[45:0] T23745;
  wire[45:0] T23746;
  wire T23747;
  wire[46:0] T23748;
  wire[46:0] T23749;
  wire T23750;
  wire T23751;
  wire T23752;
  wire T23753;
  wire T23754;
  wire T23755;
  wire T23756;
  wire T23757;
  wire[47:0] T23758;
  wire[46:0] T23759;
  wire[46:0] T23760;
  wire[46:0] T23761;
  wire[46:0] T23762;
  wire[46:0] T23763;
  wire[46:0] T23764;
  wire[46:0] T23765;
  wire[46:0] twiddle4_1_128_real;
  wire[46:0] T23766;
  wire[45:0] T23767;
  wire[45:0] T23768;
  wire T23769;
  wire[46:0] T23770;
  wire[46:0] T23771;
  wire[46:0] twiddle4_1_129_real;
  wire[46:0] T23772;
  wire[45:0] T23773;
  wire[45:0] T23774;
  wire T23775;
  wire[46:0] T23776;
  wire[46:0] T23777;
  wire T23778;
  wire[46:0] T23779;
  wire[46:0] twiddle4_1_130_real;
  wire[46:0] T23780;
  wire[45:0] T23781;
  wire[45:0] T23782;
  wire T23783;
  wire[46:0] T23784;
  wire[46:0] T23785;
  wire[46:0] twiddle4_1_131_real;
  wire[46:0] T23786;
  wire[45:0] T23787;
  wire[45:0] T23788;
  wire T23789;
  wire[46:0] T23790;
  wire[46:0] T23791;
  wire T23792;
  wire T23793;
  wire[46:0] T23794;
  wire[46:0] T23795;
  wire[46:0] twiddle4_1_132_real;
  wire[46:0] T23796;
  wire[45:0] T23797;
  wire[45:0] T23798;
  wire T23799;
  wire[46:0] T23800;
  wire[46:0] T23801;
  wire[46:0] twiddle4_1_133_real;
  wire[46:0] T23802;
  wire[45:0] T23803;
  wire[45:0] T23804;
  wire T23805;
  wire[46:0] T23806;
  wire[46:0] T23807;
  wire T23808;
  wire[46:0] T23809;
  wire[46:0] twiddle4_1_134_real;
  wire[46:0] T23810;
  wire[45:0] T23811;
  wire[45:0] T23812;
  wire T23813;
  wire[46:0] T23814;
  wire[46:0] T23815;
  wire[46:0] twiddle4_1_135_real;
  wire[46:0] T23816;
  wire[45:0] T23817;
  wire[45:0] T23818;
  wire T23819;
  wire[46:0] T23820;
  wire[46:0] T23821;
  wire T23822;
  wire T23823;
  wire T23824;
  wire[46:0] T23825;
  wire[46:0] T23826;
  wire[46:0] T23827;
  wire[46:0] twiddle4_1_136_real;
  wire[46:0] T23828;
  wire[45:0] T23829;
  wire[45:0] T23830;
  wire T23831;
  wire[46:0] T23832;
  wire[46:0] T23833;
  wire[46:0] twiddle4_1_137_real;
  wire[46:0] T23834;
  wire[45:0] T23835;
  wire[45:0] T23836;
  wire T23837;
  wire[46:0] T23838;
  wire[46:0] T23839;
  wire T23840;
  wire[46:0] T23841;
  wire[46:0] twiddle4_1_138_real;
  wire[46:0] T23842;
  wire[45:0] T23843;
  wire[45:0] T23844;
  wire T23845;
  wire[46:0] T23846;
  wire[46:0] T23847;
  wire[46:0] twiddle4_1_139_real;
  wire[46:0] T23848;
  wire[45:0] T23849;
  wire[45:0] T23850;
  wire T23851;
  wire[46:0] T23852;
  wire[46:0] T23853;
  wire T23854;
  wire T23855;
  wire[46:0] T23856;
  wire[46:0] T23857;
  wire[46:0] twiddle4_1_140_real;
  wire[46:0] T23858;
  wire[45:0] T23859;
  wire[45:0] T23860;
  wire T23861;
  wire[46:0] T23862;
  wire[46:0] T23863;
  wire[46:0] twiddle4_1_141_real;
  wire[46:0] T23864;
  wire[45:0] T23865;
  wire[45:0] T23866;
  wire T23867;
  wire[46:0] T23868;
  wire[46:0] T23869;
  wire T23870;
  wire[46:0] T23871;
  wire[46:0] twiddle4_1_142_real;
  wire[46:0] T23872;
  wire[45:0] T23873;
  wire[45:0] T23874;
  wire T23875;
  wire[46:0] T23876;
  wire[46:0] T23877;
  wire[46:0] twiddle4_1_143_real;
  wire[46:0] T23878;
  wire[45:0] T23879;
  wire[45:0] T23880;
  wire T23881;
  wire[46:0] T23882;
  wire[46:0] T23883;
  wire T23884;
  wire T23885;
  wire T23886;
  wire T23887;
  wire[46:0] T23888;
  wire[46:0] T23889;
  wire[46:0] T23890;
  wire[46:0] T23891;
  wire[46:0] twiddle4_1_144_real;
  wire[46:0] T23892;
  wire[45:0] T23893;
  wire[45:0] T23894;
  wire T23895;
  wire[46:0] T23896;
  wire[46:0] T23897;
  wire[46:0] twiddle4_1_145_real;
  wire[46:0] T23898;
  wire[45:0] T23899;
  wire[45:0] T23900;
  wire T23901;
  wire[46:0] T23902;
  wire[46:0] T23903;
  wire T23904;
  wire[46:0] T23905;
  wire[46:0] twiddle4_1_146_real;
  wire[46:0] T23906;
  wire[45:0] T23907;
  wire[45:0] T23908;
  wire T23909;
  wire[46:0] T23910;
  wire[46:0] T23911;
  wire[46:0] twiddle4_1_147_real;
  wire[46:0] T23912;
  wire[45:0] T23913;
  wire[45:0] T23914;
  wire T23915;
  wire[46:0] T23916;
  wire[46:0] T23917;
  wire T23918;
  wire T23919;
  wire[46:0] T23920;
  wire[46:0] T23921;
  wire[46:0] twiddle4_1_148_real;
  wire[46:0] T23922;
  wire[45:0] T23923;
  wire[45:0] T23924;
  wire T23925;
  wire[46:0] T23926;
  wire[46:0] T23927;
  wire[46:0] twiddle4_1_149_real;
  wire[46:0] T23928;
  wire[45:0] T23929;
  wire[45:0] T23930;
  wire T23931;
  wire[46:0] T23932;
  wire[46:0] T23933;
  wire T23934;
  wire[46:0] T23935;
  wire[46:0] twiddle4_1_150_real;
  wire[46:0] T23936;
  wire[45:0] T23937;
  wire[45:0] T23938;
  wire T23939;
  wire[46:0] T23940;
  wire[46:0] T23941;
  wire[46:0] twiddle4_1_151_real;
  wire[46:0] T23942;
  wire[45:0] T23943;
  wire[45:0] T23944;
  wire T23945;
  wire[46:0] T23946;
  wire[46:0] T23947;
  wire T23948;
  wire T23949;
  wire T23950;
  wire[46:0] T23951;
  wire[46:0] T23952;
  wire[46:0] T23953;
  wire[46:0] twiddle4_1_152_real;
  wire[46:0] T23954;
  wire[45:0] T23955;
  wire[45:0] T23956;
  wire T23957;
  wire[46:0] T23958;
  wire[46:0] T23959;
  wire[46:0] twiddle4_1_153_real;
  wire[46:0] T23960;
  wire[45:0] T23961;
  wire[45:0] T23962;
  wire T23963;
  wire[46:0] T23964;
  wire[46:0] T23965;
  wire T23966;
  wire[46:0] T23967;
  wire[46:0] twiddle4_1_154_real;
  wire[46:0] T23968;
  wire[45:0] T23969;
  wire[45:0] T23970;
  wire T23971;
  wire[46:0] T23972;
  wire[46:0] T23973;
  wire[46:0] twiddle4_1_155_real;
  wire[46:0] T23974;
  wire[45:0] T23975;
  wire[45:0] T23976;
  wire T23977;
  wire[46:0] T23978;
  wire[46:0] T23979;
  wire T23980;
  wire T23981;
  wire[46:0] T23982;
  wire[46:0] T23983;
  wire[46:0] twiddle4_1_156_real;
  wire[46:0] T23984;
  wire[45:0] T23985;
  wire[45:0] T23986;
  wire T23987;
  wire[46:0] T23988;
  wire[46:0] T23989;
  wire[46:0] twiddle4_1_157_real;
  wire[46:0] T23990;
  wire[45:0] T23991;
  wire[45:0] T23992;
  wire T23993;
  wire[46:0] T23994;
  wire[46:0] T23995;
  wire T23996;
  wire[46:0] T23997;
  wire[46:0] twiddle4_1_158_real;
  wire[46:0] T23998;
  wire[45:0] T23999;
  wire[45:0] T24000;
  wire T24001;
  wire[46:0] T24002;
  wire[46:0] T24003;
  wire[46:0] twiddle4_1_159_real;
  wire[46:0] T24004;
  wire[45:0] T24005;
  wire[45:0] T24006;
  wire T24007;
  wire[46:0] T24008;
  wire[46:0] T24009;
  wire T24010;
  wire T24011;
  wire T24012;
  wire T24013;
  wire T24014;
  wire[46:0] T24015;
  wire[46:0] T24016;
  wire[46:0] T24017;
  wire[46:0] T24018;
  wire[46:0] T24019;
  wire[46:0] twiddle4_1_160_real;
  wire[46:0] T24020;
  wire[45:0] T24021;
  wire[45:0] T24022;
  wire T24023;
  wire[46:0] T24024;
  wire[46:0] T24025;
  wire[46:0] twiddle4_1_161_real;
  wire[46:0] T24026;
  wire[45:0] T24027;
  wire[45:0] T24028;
  wire T24029;
  wire[46:0] T24030;
  wire[46:0] T24031;
  wire T24032;
  wire[46:0] T24033;
  wire[46:0] twiddle4_1_162_real;
  wire[46:0] T24034;
  wire[45:0] T24035;
  wire[45:0] T24036;
  wire T24037;
  wire[46:0] T24038;
  wire[46:0] T24039;
  wire[46:0] twiddle4_1_163_real;
  wire[46:0] T24040;
  wire[45:0] T24041;
  wire[45:0] T24042;
  wire T24043;
  wire[46:0] T24044;
  wire[46:0] T24045;
  wire T24046;
  wire T24047;
  wire[46:0] T24048;
  wire[46:0] T24049;
  wire[46:0] twiddle4_1_164_real;
  wire[46:0] T24050;
  wire[45:0] T24051;
  wire[45:0] T24052;
  wire T24053;
  wire[46:0] T24054;
  wire[46:0] T24055;
  wire[46:0] twiddle4_1_165_real;
  wire[46:0] T24056;
  wire[45:0] T24057;
  wire[45:0] T24058;
  wire T24059;
  wire[46:0] T24060;
  wire[46:0] T24061;
  wire T24062;
  wire[46:0] T24063;
  wire[46:0] twiddle4_1_166_real;
  wire[46:0] T24064;
  wire[45:0] T24065;
  wire[45:0] T24066;
  wire T24067;
  wire[46:0] T24068;
  wire[46:0] T24069;
  wire[46:0] twiddle4_1_167_real;
  wire[46:0] T24070;
  wire[45:0] T24071;
  wire[45:0] T24072;
  wire T24073;
  wire[46:0] T24074;
  wire[46:0] T24075;
  wire T24076;
  wire T24077;
  wire T24078;
  wire[46:0] T24079;
  wire[46:0] T24080;
  wire[46:0] T24081;
  wire[46:0] twiddle4_1_168_real;
  wire[46:0] T24082;
  wire[45:0] T24083;
  wire[45:0] T24084;
  wire T24085;
  wire[46:0] T24086;
  wire[46:0] T24087;
  wire[46:0] twiddle4_1_169_real;
  wire[46:0] T24088;
  wire[45:0] T24089;
  wire[45:0] T24090;
  wire T24091;
  wire[46:0] T24092;
  wire[46:0] T24093;
  wire T24094;
  wire[46:0] T24095;
  wire[46:0] twiddle4_1_170_real;
  wire[46:0] T24096;
  wire[45:0] T24097;
  wire[45:0] T24098;
  wire T24099;
  wire[46:0] T24100;
  wire[46:0] T24101;
  wire[46:0] twiddle4_1_171_real;
  wire[46:0] T24102;
  wire[46:0] T24103;
  wire[46:0] T24104;
  wire[46:0] T24105;
  wire T24106;
  wire T24107;
  wire[46:0] T24108;
  wire[46:0] T24109;
  wire[46:0] twiddle4_1_172_real;
  wire[46:0] T24110;
  wire[46:0] T24111;
  wire[46:0] T24112;
  wire[46:0] T24113;
  wire[46:0] twiddle4_1_173_real;
  wire[46:0] T24114;
  wire[46:0] T24115;
  wire[46:0] T24116;
  wire[46:0] T24117;
  wire T24118;
  wire[46:0] T24119;
  wire[46:0] twiddle4_1_174_real;
  wire[46:0] T24120;
  wire[46:0] T24121;
  wire[46:0] T24122;
  wire[46:0] T24123;
  wire[46:0] twiddle4_1_175_real;
  wire[46:0] T24124;
  wire[46:0] T24125;
  wire[46:0] T24126;
  wire[46:0] T24127;
  wire T24128;
  wire T24129;
  wire T24130;
  wire T24131;
  wire[46:0] T24132;
  wire[46:0] T24133;
  wire[46:0] T24134;
  wire[46:0] T24135;
  wire[46:0] twiddle4_1_176_real;
  wire[46:0] T24136;
  wire[46:0] T24137;
  wire[46:0] T24138;
  wire[46:0] T24139;
  wire[46:0] twiddle4_1_177_real;
  wire[46:0] T24140;
  wire[46:0] T24141;
  wire[46:0] T24142;
  wire[46:0] T24143;
  wire T24144;
  wire[46:0] T24145;
  wire[46:0] twiddle4_1_178_real;
  wire[46:0] T24146;
  wire[46:0] T24147;
  wire[46:0] T24148;
  wire[46:0] T24149;
  wire[46:0] twiddle4_1_179_real;
  wire[46:0] T24150;
  wire[46:0] T24151;
  wire[46:0] T24152;
  wire[46:0] T24153;
  wire T24154;
  wire T24155;
  wire[46:0] T24156;
  wire[46:0] T24157;
  wire[46:0] twiddle4_1_180_real;
  wire[46:0] T24158;
  wire[46:0] T24159;
  wire[46:0] T24160;
  wire[46:0] T24161;
  wire[46:0] twiddle4_1_181_real;
  wire[46:0] T24162;
  wire[46:0] T24163;
  wire[46:0] T24164;
  wire[46:0] T24165;
  wire T24166;
  wire[46:0] T24167;
  wire[46:0] twiddle4_1_182_real;
  wire[46:0] T24168;
  wire[46:0] T24169;
  wire[46:0] T24170;
  wire[46:0] T24171;
  wire[46:0] twiddle4_1_183_real;
  wire[46:0] T24172;
  wire[46:0] T24173;
  wire[46:0] T24174;
  wire[46:0] T24175;
  wire T24176;
  wire T24177;
  wire T24178;
  wire[46:0] T24179;
  wire[46:0] T24180;
  wire[46:0] T24181;
  wire[46:0] twiddle4_1_184_real;
  wire[46:0] T24182;
  wire[46:0] T24183;
  wire[46:0] T24184;
  wire[46:0] T24185;
  wire[46:0] twiddle4_1_185_real;
  wire[46:0] T24186;
  wire[46:0] T24187;
  wire[46:0] T24188;
  wire[46:0] T24189;
  wire T24190;
  wire[46:0] T24191;
  wire[46:0] twiddle4_1_186_real;
  wire[46:0] T24192;
  wire[46:0] T24193;
  wire[46:0] T24194;
  wire[46:0] T24195;
  wire[46:0] twiddle4_1_187_real;
  wire[46:0] T24196;
  wire[46:0] T24197;
  wire[46:0] T24198;
  wire[46:0] T24199;
  wire T24200;
  wire T24201;
  wire[46:0] T24202;
  wire[46:0] T24203;
  wire[46:0] twiddle4_1_188_real;
  wire[46:0] T24204;
  wire[46:0] T24205;
  wire[46:0] T24206;
  wire[46:0] T24207;
  wire[46:0] twiddle4_1_189_real;
  wire[46:0] T24208;
  wire[46:0] T24209;
  wire[46:0] T24210;
  wire[46:0] T24211;
  wire T24212;
  wire[46:0] T24213;
  wire[46:0] twiddle4_1_190_real;
  wire[46:0] T24214;
  wire[46:0] T24215;
  wire[46:0] T24216;
  wire[46:0] T24217;
  wire[46:0] twiddle4_1_191_real;
  wire[46:0] T24218;
  wire[46:0] T24219;
  wire[46:0] T24220;
  wire[46:0] T24221;
  wire T24222;
  wire T24223;
  wire T24224;
  wire T24225;
  wire T24226;
  wire T24227;
  wire[46:0] T24228;
  wire[46:0] T24229;
  wire[46:0] T24230;
  wire[46:0] T24231;
  wire[46:0] T24232;
  wire[46:0] T24233;
  wire[46:0] twiddle4_1_192_real;
  wire[46:0] T24234;
  wire[46:0] T24235;
  wire[46:0] T24236;
  wire[46:0] T24237;
  wire[46:0] twiddle4_1_193_real;
  wire[46:0] T24238;
  wire[46:0] T24239;
  wire[46:0] T24240;
  wire[46:0] T24241;
  wire T24242;
  wire[46:0] T24243;
  wire[46:0] twiddle4_1_194_real;
  wire[46:0] T24244;
  wire[46:0] T24245;
  wire[46:0] T24246;
  wire[46:0] T24247;
  wire[46:0] twiddle4_1_195_real;
  wire[46:0] T24248;
  wire[46:0] T24249;
  wire[46:0] T24250;
  wire[46:0] T24251;
  wire T24252;
  wire T24253;
  wire[46:0] T24254;
  wire[46:0] T24255;
  wire[46:0] twiddle4_1_196_real;
  wire[46:0] T24256;
  wire[46:0] T24257;
  wire[46:0] T24258;
  wire[46:0] T24259;
  wire[46:0] twiddle4_1_197_real;
  wire[46:0] T24260;
  wire[46:0] T24261;
  wire[46:0] T24262;
  wire[46:0] T24263;
  wire T24264;
  wire[46:0] T24265;
  wire[46:0] twiddle4_1_198_real;
  wire[46:0] T24266;
  wire[46:0] T24267;
  wire[46:0] T24268;
  wire[46:0] T24269;
  wire[46:0] twiddle4_1_199_real;
  wire[46:0] T24270;
  wire[46:0] T24271;
  wire[46:0] T24272;
  wire[46:0] T24273;
  wire T24274;
  wire T24275;
  wire T24276;
  wire[46:0] T24277;
  wire[46:0] T24278;
  wire[46:0] T24279;
  wire[46:0] twiddle4_1_200_real;
  wire[46:0] T24280;
  wire[46:0] T24281;
  wire[46:0] T24282;
  wire[46:0] T24283;
  wire[46:0] twiddle4_1_201_real;
  wire[46:0] T24284;
  wire[46:0] T24285;
  wire[46:0] T24286;
  wire[46:0] T24287;
  wire T24288;
  wire[46:0] T24289;
  wire[46:0] twiddle4_1_202_real;
  wire[46:0] T24290;
  wire[46:0] T24291;
  wire[46:0] T24292;
  wire[46:0] T24293;
  wire[46:0] twiddle4_1_203_real;
  wire[46:0] T24294;
  wire[46:0] T24295;
  wire[46:0] T24296;
  wire[46:0] T24297;
  wire T24298;
  wire T24299;
  wire[46:0] T24300;
  wire[46:0] T24301;
  wire[46:0] twiddle4_1_204_real;
  wire[46:0] T24302;
  wire[46:0] T24303;
  wire[46:0] T24304;
  wire[46:0] T24305;
  wire[46:0] twiddle4_1_205_real;
  wire[46:0] T24306;
  wire[46:0] T24307;
  wire[46:0] T24308;
  wire[46:0] T24309;
  wire T24310;
  wire[46:0] T24311;
  wire[46:0] twiddle4_1_206_real;
  wire[46:0] T24312;
  wire[46:0] T24313;
  wire[46:0] T24314;
  wire[46:0] T24315;
  wire[46:0] twiddle4_1_207_real;
  wire[46:0] T24316;
  wire[46:0] T24317;
  wire[46:0] T24318;
  wire[46:0] T24319;
  wire T24320;
  wire T24321;
  wire T24322;
  wire T24323;
  wire[46:0] T24324;
  wire[46:0] T24325;
  wire[46:0] T24326;
  wire[46:0] T24327;
  wire[46:0] twiddle4_1_208_real;
  wire[46:0] T24328;
  wire[46:0] T24329;
  wire[46:0] T24330;
  wire[46:0] T24331;
  wire[46:0] twiddle4_1_209_real;
  wire[46:0] T24332;
  wire[46:0] T24333;
  wire[46:0] T24334;
  wire[46:0] T24335;
  wire T24336;
  wire[46:0] T24337;
  wire[46:0] twiddle4_1_210_real;
  wire[46:0] T24338;
  wire[46:0] T24339;
  wire[46:0] T24340;
  wire[46:0] T24341;
  wire[46:0] twiddle4_1_211_real;
  wire[46:0] T24342;
  wire[46:0] T24343;
  wire[46:0] T24344;
  wire[46:0] T24345;
  wire T24346;
  wire T24347;
  wire[46:0] T24348;
  wire[46:0] T24349;
  wire[46:0] twiddle4_1_212_real;
  wire[46:0] T24350;
  wire[46:0] T24351;
  wire[46:0] T24352;
  wire[46:0] T24353;
  wire[46:0] twiddle4_1_213_real;
  wire[46:0] T24354;
  wire[46:0] T24355;
  wire[46:0] T24356;
  wire[46:0] T24357;
  wire T24358;
  wire[46:0] T24359;
  wire[46:0] twiddle4_1_214_real;
  wire[46:0] T24360;
  wire[46:0] T24361;
  wire[46:0] T24362;
  wire[46:0] T24363;
  wire[46:0] twiddle4_1_215_real;
  wire[46:0] T24364;
  wire[46:0] T24365;
  wire[46:0] T24366;
  wire[46:0] T24367;
  wire T24368;
  wire T24369;
  wire T24370;
  wire[46:0] T24371;
  wire[46:0] T24372;
  wire[46:0] T24373;
  wire[46:0] twiddle4_1_216_real;
  wire[46:0] T24374;
  wire[46:0] T24375;
  wire[46:0] T24376;
  wire[46:0] T24377;
  wire[46:0] twiddle4_1_217_real;
  wire[46:0] T24378;
  wire[46:0] T24379;
  wire[46:0] T24380;
  wire[46:0] T24381;
  wire T24382;
  wire[46:0] T24383;
  wire[46:0] twiddle4_1_218_real;
  wire[46:0] T24384;
  wire[46:0] T24385;
  wire[46:0] T24386;
  wire[46:0] T24387;
  wire[46:0] twiddle4_1_219_real;
  wire[46:0] T24388;
  wire[46:0] T24389;
  wire[46:0] T24390;
  wire[46:0] T24391;
  wire T24392;
  wire T24393;
  wire[46:0] T24394;
  wire[46:0] T24395;
  wire[46:0] twiddle4_1_220_real;
  wire[46:0] T24396;
  wire[46:0] T24397;
  wire[46:0] T24398;
  wire[46:0] T24399;
  wire[46:0] twiddle4_1_221_real;
  wire[46:0] T24400;
  wire[46:0] T24401;
  wire[46:0] T24402;
  wire[46:0] T24403;
  wire T24404;
  wire[46:0] T24405;
  wire[46:0] twiddle4_1_222_real;
  wire[46:0] T24406;
  wire[46:0] T24407;
  wire[46:0] T24408;
  wire[46:0] T24409;
  wire[46:0] twiddle4_1_223_real;
  wire[46:0] T24410;
  wire[46:0] T24411;
  wire[46:0] T24412;
  wire[46:0] T24413;
  wire T24414;
  wire T24415;
  wire T24416;
  wire T24417;
  wire T24418;
  wire[46:0] T24419;
  wire[46:0] T24420;
  wire[46:0] T24421;
  wire[46:0] T24422;
  wire[46:0] T24423;
  wire[46:0] twiddle4_1_224_real;
  wire[46:0] T24424;
  wire[46:0] T24425;
  wire[46:0] T24426;
  wire[46:0] T24427;
  wire[46:0] twiddle4_1_225_real;
  wire[46:0] T24428;
  wire[46:0] T24429;
  wire[46:0] T24430;
  wire[46:0] T24431;
  wire T24432;
  wire[46:0] T24433;
  wire[46:0] twiddle4_1_226_real;
  wire[46:0] T24434;
  wire[46:0] T24435;
  wire[46:0] T24436;
  wire[46:0] T24437;
  wire[46:0] twiddle4_1_227_real;
  wire[46:0] T24438;
  wire[46:0] T24439;
  wire[46:0] T24440;
  wire[46:0] T24441;
  wire T24442;
  wire T24443;
  wire[46:0] T24444;
  wire[46:0] T24445;
  wire[46:0] twiddle4_1_228_real;
  wire[46:0] T24446;
  wire[46:0] T24447;
  wire[46:0] T24448;
  wire[46:0] T24449;
  wire[46:0] twiddle4_1_229_real;
  wire[46:0] T24450;
  wire[46:0] T24451;
  wire[46:0] T24452;
  wire[46:0] T24453;
  wire T24454;
  wire[46:0] T24455;
  wire[46:0] twiddle4_1_230_real;
  wire[46:0] T24456;
  wire[46:0] T24457;
  wire[46:0] T24458;
  wire[46:0] T24459;
  wire[46:0] twiddle4_1_231_real;
  wire[46:0] T24460;
  wire[46:0] T24461;
  wire[46:0] T24462;
  wire[46:0] T24463;
  wire T24464;
  wire T24465;
  wire T24466;
  wire[46:0] T24467;
  wire[46:0] T24468;
  wire[46:0] T24469;
  wire[46:0] twiddle4_1_232_real;
  wire[46:0] T24470;
  wire[46:0] T24471;
  wire[46:0] T24472;
  wire[46:0] T24473;
  wire[46:0] twiddle4_1_233_real;
  wire[46:0] T24474;
  wire[46:0] T24475;
  wire[46:0] T24476;
  wire[46:0] T24477;
  wire T24478;
  wire[46:0] T24479;
  wire[46:0] twiddle4_1_234_real;
  wire[46:0] T24480;
  wire[46:0] T24481;
  wire[46:0] T24482;
  wire[46:0] T24483;
  wire[46:0] twiddle4_1_235_real;
  wire[46:0] T24484;
  wire[46:0] T24485;
  wire[46:0] T24486;
  wire[46:0] T24487;
  wire T24488;
  wire T24489;
  wire[46:0] T24490;
  wire[46:0] T24491;
  wire[46:0] twiddle4_1_236_real;
  wire[46:0] T24492;
  wire[46:0] T24493;
  wire[46:0] T24494;
  wire[46:0] T24495;
  wire[46:0] twiddle4_1_237_real;
  wire[46:0] T24496;
  wire[46:0] T24497;
  wire[46:0] T24498;
  wire[46:0] T24499;
  wire T24500;
  wire[46:0] T24501;
  wire[46:0] twiddle4_1_238_real;
  wire[46:0] T24502;
  wire[46:0] T24503;
  wire[46:0] T24504;
  wire[46:0] T24505;
  wire[46:0] twiddle4_1_239_real;
  wire[46:0] T24506;
  wire[46:0] T24507;
  wire[46:0] T24508;
  wire[46:0] T24509;
  wire T24510;
  wire T24511;
  wire T24512;
  wire T24513;
  wire[46:0] T24514;
  wire[46:0] T24515;
  wire[46:0] T24516;
  wire[46:0] T24517;
  wire[46:0] twiddle4_1_240_real;
  wire[46:0] T24518;
  wire[46:0] T24519;
  wire[46:0] T24520;
  wire[46:0] T24521;
  wire[46:0] twiddle4_1_241_real;
  wire[46:0] T24522;
  wire[46:0] T24523;
  wire[46:0] T24524;
  wire[46:0] T24525;
  wire T24526;
  wire[46:0] T24527;
  wire[46:0] twiddle4_1_242_real;
  wire[46:0] T24528;
  wire[46:0] T24529;
  wire[46:0] T24530;
  wire[46:0] T24531;
  wire[46:0] twiddle4_1_243_real;
  wire[46:0] T24532;
  wire[46:0] T24533;
  wire[46:0] T24534;
  wire[46:0] T24535;
  wire T24536;
  wire T24537;
  wire[46:0] T24538;
  wire[46:0] T24539;
  wire[46:0] twiddle4_1_244_real;
  wire[46:0] T24540;
  wire[46:0] T24541;
  wire[46:0] T24542;
  wire[46:0] T24543;
  wire[46:0] twiddle4_1_245_real;
  wire[46:0] T24544;
  wire[46:0] T24545;
  wire[46:0] T24546;
  wire[46:0] T24547;
  wire T24548;
  wire[46:0] T24549;
  wire[46:0] twiddle4_1_246_real;
  wire[46:0] T24550;
  wire[46:0] T24551;
  wire[46:0] T24552;
  wire[46:0] T24553;
  wire[46:0] twiddle4_1_247_real;
  wire[46:0] T24554;
  wire[46:0] T24555;
  wire[46:0] T24556;
  wire[46:0] T24557;
  wire T24558;
  wire T24559;
  wire T24560;
  wire[46:0] T24561;
  wire[46:0] T24562;
  wire[46:0] T24563;
  wire[46:0] twiddle4_1_248_real;
  wire[46:0] T24564;
  wire[46:0] T24565;
  wire[46:0] T24566;
  wire[46:0] T24567;
  wire[46:0] twiddle4_1_249_real;
  wire[46:0] T24568;
  wire[46:0] T24569;
  wire[46:0] T24570;
  wire[46:0] T24571;
  wire T24572;
  wire[46:0] T24573;
  wire[46:0] twiddle4_1_250_real;
  wire[46:0] T24574;
  wire[46:0] T24575;
  wire[46:0] T24576;
  wire[46:0] T24577;
  wire[46:0] twiddle4_1_251_real;
  wire[46:0] T24578;
  wire[46:0] T24579;
  wire[46:0] T24580;
  wire[46:0] T24581;
  wire T24582;
  wire T24583;
  wire[46:0] T24584;
  wire[46:0] T24585;
  wire[46:0] twiddle4_1_252_real;
  wire[46:0] T24586;
  wire[46:0] T24587;
  wire[46:0] T24588;
  wire[46:0] T24589;
  wire[46:0] twiddle4_1_253_real;
  wire[46:0] T24590;
  wire[46:0] T24591;
  wire[46:0] T24592;
  wire[46:0] T24593;
  wire T24594;
  wire[46:0] T24595;
  wire[46:0] twiddle4_1_254_real;
  wire[46:0] T24596;
  wire[46:0] T24597;
  wire[46:0] T24598;
  wire[46:0] T24599;
  wire[46:0] twiddle4_1_255_real;
  wire[46:0] T24600;
  wire[46:0] T24601;
  wire[46:0] T24602;
  wire[46:0] T24603;
  wire T24604;
  wire T24605;
  wire T24606;
  wire T24607;
  wire T24608;
  wire T24609;
  wire T24610;
  wire T24611;
  wire T24612;
  wire[47:0] T24613;
  wire[46:0] T24614;
  wire[46:0] T24615;
  wire[46:0] T24616;
  wire[46:0] T24617;
  wire[46:0] T24618;
  wire[46:0] T24619;
  wire[46:0] T24620;
  wire[46:0] T24621;
  wire[46:0] twiddle4_1_256_real;
  wire[46:0] T24622;
  wire[46:0] T24623;
  wire[46:0] T24624;
  wire[46:0] T24625;
  wire[46:0] twiddle4_1_257_real;
  wire[46:0] T24626;
  wire[46:0] T24627;
  wire[46:0] T24628;
  wire[46:0] T24629;
  wire T24630;
  wire[46:0] T24631;
  wire[46:0] twiddle4_1_258_real;
  wire[46:0] T24632;
  wire[46:0] T24633;
  wire[46:0] T24634;
  wire[46:0] T24635;
  wire[46:0] twiddle4_1_259_real;
  wire[46:0] T24636;
  wire[46:0] T24637;
  wire[46:0] T24638;
  wire[46:0] T24639;
  wire T24640;
  wire T24641;
  wire[46:0] T24642;
  wire[46:0] T24643;
  wire[46:0] twiddle4_1_260_real;
  wire[46:0] T24644;
  wire[46:0] T24645;
  wire[46:0] T24646;
  wire[46:0] T24647;
  wire[46:0] twiddle4_1_261_real;
  wire[46:0] T24648;
  wire[46:0] T24649;
  wire[46:0] T24650;
  wire[46:0] T24651;
  wire T24652;
  wire[46:0] T24653;
  wire[46:0] twiddle4_1_262_real;
  wire[46:0] T24654;
  wire[46:0] T24655;
  wire[46:0] T24656;
  wire[46:0] T24657;
  wire[46:0] twiddle4_1_263_real;
  wire[46:0] T24658;
  wire[46:0] T24659;
  wire[46:0] T24660;
  wire[46:0] T24661;
  wire T24662;
  wire T24663;
  wire T24664;
  wire[46:0] T24665;
  wire[46:0] T24666;
  wire[46:0] T24667;
  wire[46:0] twiddle4_1_264_real;
  wire[46:0] T24668;
  wire[46:0] T24669;
  wire[46:0] T24670;
  wire[46:0] T24671;
  wire[46:0] twiddle4_1_265_real;
  wire[46:0] T24672;
  wire[46:0] T24673;
  wire[46:0] T24674;
  wire[46:0] T24675;
  wire T24676;
  wire[46:0] T24677;
  wire[46:0] twiddle4_1_266_real;
  wire[46:0] T24678;
  wire[46:0] T24679;
  wire[46:0] T24680;
  wire[46:0] T24681;
  wire[46:0] twiddle4_1_267_real;
  wire[46:0] T24682;
  wire[46:0] T24683;
  wire[46:0] T24684;
  wire[46:0] T24685;
  wire T24686;
  wire T24687;
  wire[46:0] T24688;
  wire[46:0] T24689;
  wire[46:0] twiddle4_1_268_real;
  wire[46:0] T24690;
  wire[46:0] T24691;
  wire[46:0] T24692;
  wire[46:0] T24693;
  wire[46:0] twiddle4_1_269_real;
  wire[46:0] T24694;
  wire[46:0] T24695;
  wire[46:0] T24696;
  wire[46:0] T24697;
  wire T24698;
  wire[46:0] T24699;
  wire[46:0] twiddle4_1_270_real;
  wire[46:0] T24700;
  wire[46:0] T24701;
  wire[46:0] T24702;
  wire[46:0] T24703;
  wire[46:0] twiddle4_1_271_real;
  wire[46:0] T24704;
  wire[46:0] T24705;
  wire[46:0] T24706;
  wire[46:0] T24707;
  wire T24708;
  wire T24709;
  wire T24710;
  wire T24711;
  wire[46:0] T24712;
  wire[46:0] T24713;
  wire[46:0] T24714;
  wire[46:0] T24715;
  wire[46:0] twiddle4_1_272_real;
  wire[46:0] T24716;
  wire[46:0] T24717;
  wire[46:0] T24718;
  wire[46:0] T24719;
  wire[46:0] twiddle4_1_273_real;
  wire[46:0] T24720;
  wire[46:0] T24721;
  wire[46:0] T24722;
  wire[46:0] T24723;
  wire T24724;
  wire[46:0] T24725;
  wire[46:0] twiddle4_1_274_real;
  wire[46:0] T24726;
  wire[46:0] T24727;
  wire[46:0] T24728;
  wire[46:0] T24729;
  wire[46:0] twiddle4_1_275_real;
  wire[46:0] T24730;
  wire[46:0] T24731;
  wire[46:0] T24732;
  wire[46:0] T24733;
  wire T24734;
  wire T24735;
  wire[46:0] T24736;
  wire[46:0] T24737;
  wire[46:0] twiddle4_1_276_real;
  wire[46:0] T24738;
  wire[46:0] T24739;
  wire[46:0] T24740;
  wire[46:0] T24741;
  wire[46:0] twiddle4_1_277_real;
  wire[46:0] T24742;
  wire[46:0] T24743;
  wire[46:0] T24744;
  wire[46:0] T24745;
  wire T24746;
  wire[46:0] T24747;
  wire[46:0] twiddle4_1_278_real;
  wire[46:0] T24748;
  wire[46:0] T24749;
  wire[46:0] T24750;
  wire[46:0] T24751;
  wire[46:0] twiddle4_1_279_real;
  wire[46:0] T24752;
  wire[46:0] T24753;
  wire[46:0] T24754;
  wire[46:0] T24755;
  wire T24756;
  wire T24757;
  wire T24758;
  wire[46:0] T24759;
  wire[46:0] T24760;
  wire[46:0] T24761;
  wire[46:0] twiddle4_1_280_real;
  wire[46:0] T24762;
  wire[46:0] T24763;
  wire[46:0] T24764;
  wire[46:0] T24765;
  wire[46:0] twiddle4_1_281_real;
  wire[46:0] T24766;
  wire[46:0] T24767;
  wire[46:0] T24768;
  wire[46:0] T24769;
  wire T24770;
  wire[46:0] T24771;
  wire[46:0] twiddle4_1_282_real;
  wire[46:0] T24772;
  wire[46:0] T24773;
  wire[46:0] T24774;
  wire[46:0] T24775;
  wire[46:0] twiddle4_1_283_real;
  wire[46:0] T24776;
  wire[46:0] T24777;
  wire[46:0] T24778;
  wire[46:0] T24779;
  wire T24780;
  wire T24781;
  wire[46:0] T24782;
  wire[46:0] T24783;
  wire[46:0] twiddle4_1_284_real;
  wire[46:0] T24784;
  wire[46:0] T24785;
  wire[46:0] T24786;
  wire[46:0] T24787;
  wire[46:0] twiddle4_1_285_real;
  wire[46:0] T24788;
  wire[46:0] T24789;
  wire[46:0] T24790;
  wire[46:0] T24791;
  wire T24792;
  wire[46:0] T24793;
  wire[46:0] twiddle4_1_286_real;
  wire[46:0] T24794;
  wire[46:0] T24795;
  wire[46:0] T24796;
  wire[46:0] T24797;
  wire[46:0] twiddle4_1_287_real;
  wire[46:0] T24798;
  wire[46:0] T24799;
  wire[46:0] T24800;
  wire[46:0] T24801;
  wire T24802;
  wire T24803;
  wire T24804;
  wire T24805;
  wire T24806;
  wire[46:0] T24807;
  wire[46:0] T24808;
  wire[46:0] T24809;
  wire[46:0] T24810;
  wire[46:0] T24811;
  wire[46:0] twiddle4_1_288_real;
  wire[46:0] T24812;
  wire[46:0] T24813;
  wire[46:0] T24814;
  wire[46:0] T24815;
  wire[46:0] twiddle4_1_289_real;
  wire[46:0] T24816;
  wire[46:0] T24817;
  wire[46:0] T24818;
  wire[46:0] T24819;
  wire T24820;
  wire[46:0] T24821;
  wire[46:0] twiddle4_1_290_real;
  wire[46:0] T24822;
  wire[46:0] T24823;
  wire[46:0] T24824;
  wire[46:0] T24825;
  wire[46:0] twiddle4_1_291_real;
  wire[46:0] T24826;
  wire[46:0] T24827;
  wire[46:0] T24828;
  wire[46:0] T24829;
  wire T24830;
  wire T24831;
  wire[46:0] T24832;
  wire[46:0] T24833;
  wire[46:0] twiddle4_1_292_real;
  wire[46:0] T24834;
  wire[46:0] T24835;
  wire[46:0] T24836;
  wire[46:0] T24837;
  wire[46:0] twiddle4_1_293_real;
  wire[46:0] T24838;
  wire[46:0] T24839;
  wire[46:0] T24840;
  wire[46:0] T24841;
  wire T24842;
  wire[46:0] T24843;
  wire[46:0] twiddle4_1_294_real;
  wire[46:0] T24844;
  wire[46:0] T24845;
  wire[46:0] T24846;
  wire[46:0] T24847;
  wire[46:0] twiddle4_1_295_real;
  wire[46:0] T24848;
  wire[46:0] T24849;
  wire[46:0] T24850;
  wire[46:0] T24851;
  wire T24852;
  wire T24853;
  wire T24854;
  wire[46:0] T24855;
  wire[46:0] T24856;
  wire[46:0] T24857;
  wire[46:0] twiddle4_1_296_real;
  wire[46:0] T24858;
  wire[46:0] T24859;
  wire[46:0] T24860;
  wire[46:0] T24861;
  wire[46:0] twiddle4_1_297_real;
  wire[46:0] T24862;
  wire[46:0] T24863;
  wire[46:0] T24864;
  wire[46:0] T24865;
  wire T24866;
  wire[46:0] T24867;
  wire[46:0] twiddle4_1_298_real;
  wire[46:0] T24868;
  wire[46:0] T24869;
  wire[46:0] T24870;
  wire[46:0] T24871;
  wire[46:0] twiddle4_1_299_real;
  wire[46:0] T24872;
  wire[46:0] T24873;
  wire[46:0] T24874;
  wire[46:0] T24875;
  wire T24876;
  wire T24877;
  wire[46:0] T24878;
  wire[46:0] T24879;
  wire[46:0] twiddle4_1_300_real;
  wire[46:0] T24880;
  wire[46:0] T24881;
  wire[46:0] T24882;
  wire[46:0] T24883;
  wire[46:0] twiddle4_1_301_real;
  wire[46:0] T24884;
  wire[46:0] T24885;
  wire[46:0] T24886;
  wire[46:0] T24887;
  wire T24888;
  wire[46:0] T24889;
  wire[46:0] twiddle4_1_302_real;
  wire[46:0] T24890;
  wire[46:0] T24891;
  wire[46:0] T24892;
  wire[46:0] T24893;
  wire[46:0] twiddle4_1_303_real;
  wire[46:0] T24894;
  wire[46:0] T24895;
  wire[46:0] T24896;
  wire[46:0] T24897;
  wire T24898;
  wire T24899;
  wire T24900;
  wire T24901;
  wire[46:0] T24902;
  wire[46:0] T24903;
  wire[46:0] T24904;
  wire[46:0] T24905;
  wire[46:0] twiddle4_1_304_real;
  wire[46:0] T24906;
  wire[46:0] T24907;
  wire[46:0] T24908;
  wire[46:0] T24909;
  wire[46:0] twiddle4_1_305_real;
  wire[46:0] T24910;
  wire[46:0] T24911;
  wire[46:0] T24912;
  wire[46:0] T24913;
  wire T24914;
  wire[46:0] T24915;
  wire[46:0] twiddle4_1_306_real;
  wire[46:0] T24916;
  wire[46:0] T24917;
  wire[46:0] T24918;
  wire[46:0] T24919;
  wire[46:0] twiddle4_1_307_real;
  wire[46:0] T24920;
  wire[46:0] T24921;
  wire[46:0] T24922;
  wire[46:0] T24923;
  wire T24924;
  wire T24925;
  wire[46:0] T24926;
  wire[46:0] T24927;
  wire[46:0] twiddle4_1_308_real;
  wire[46:0] T24928;
  wire[46:0] T24929;
  wire[46:0] T24930;
  wire[46:0] T24931;
  wire[46:0] twiddle4_1_309_real;
  wire[46:0] T24932;
  wire[46:0] T24933;
  wire[46:0] T24934;
  wire[46:0] T24935;
  wire T24936;
  wire[46:0] T24937;
  wire[46:0] twiddle4_1_310_real;
  wire[46:0] T24938;
  wire[46:0] T24939;
  wire[46:0] T24940;
  wire[46:0] T24941;
  wire[46:0] twiddle4_1_311_real;
  wire[46:0] T24942;
  wire[46:0] T24943;
  wire[46:0] T24944;
  wire[46:0] T24945;
  wire T24946;
  wire T24947;
  wire T24948;
  wire[46:0] T24949;
  wire[46:0] T24950;
  wire[46:0] T24951;
  wire[46:0] twiddle4_1_312_real;
  wire[46:0] T24952;
  wire[46:0] T24953;
  wire[46:0] T24954;
  wire[46:0] T24955;
  wire[46:0] twiddle4_1_313_real;
  wire[46:0] T24956;
  wire[46:0] T24957;
  wire[46:0] T24958;
  wire[46:0] T24959;
  wire T24960;
  wire[46:0] T24961;
  wire[46:0] twiddle4_1_314_real;
  wire[46:0] T24962;
  wire[46:0] T24963;
  wire[46:0] T24964;
  wire[46:0] T24965;
  wire[46:0] twiddle4_1_315_real;
  wire[46:0] T24966;
  wire[46:0] T24967;
  wire[46:0] T24968;
  wire[46:0] T24969;
  wire T24970;
  wire T24971;
  wire[46:0] T24972;
  wire[46:0] T24973;
  wire[46:0] twiddle4_1_316_real;
  wire[46:0] T24974;
  wire[46:0] T24975;
  wire[46:0] T24976;
  wire[46:0] T24977;
  wire[46:0] twiddle4_1_317_real;
  wire[46:0] T24978;
  wire[46:0] T24979;
  wire[46:0] T24980;
  wire[46:0] T24981;
  wire T24982;
  wire[46:0] T24983;
  wire[46:0] twiddle4_1_318_real;
  wire[46:0] T24984;
  wire[46:0] T24985;
  wire[46:0] T24986;
  wire[46:0] T24987;
  wire[46:0] twiddle4_1_319_real;
  wire[46:0] T24988;
  wire[46:0] T24989;
  wire[46:0] T24990;
  wire[46:0] T24991;
  wire T24992;
  wire T24993;
  wire T24994;
  wire T24995;
  wire T24996;
  wire T24997;
  wire[46:0] T24998;
  wire[46:0] T24999;
  wire[46:0] T25000;
  wire[46:0] T25001;
  wire[46:0] T25002;
  wire[46:0] T25003;
  wire[46:0] twiddle4_1_320_real;
  wire[46:0] T25004;
  wire[46:0] T25005;
  wire[46:0] T25006;
  wire[46:0] T25007;
  wire[46:0] twiddle4_1_321_real;
  wire[46:0] T25008;
  wire[46:0] T25009;
  wire[46:0] T25010;
  wire[46:0] T25011;
  wire T25012;
  wire[46:0] T25013;
  wire[46:0] twiddle4_1_322_real;
  wire[46:0] T25014;
  wire[46:0] T25015;
  wire[46:0] T25016;
  wire[46:0] T25017;
  wire[46:0] twiddle4_1_323_real;
  wire[46:0] T25018;
  wire[46:0] T25019;
  wire[46:0] T25020;
  wire[46:0] T25021;
  wire T25022;
  wire T25023;
  wire[46:0] T25024;
  wire[46:0] T25025;
  wire[46:0] twiddle4_1_324_real;
  wire[46:0] T25026;
  wire[46:0] T25027;
  wire[46:0] T25028;
  wire[46:0] T25029;
  wire[46:0] twiddle4_1_325_real;
  wire[46:0] T25030;
  wire[46:0] T25031;
  wire[46:0] T25032;
  wire[46:0] T25033;
  wire T25034;
  wire[46:0] T25035;
  wire[46:0] twiddle4_1_326_real;
  wire[46:0] T25036;
  wire[46:0] T25037;
  wire[46:0] T25038;
  wire[46:0] T25039;
  wire[46:0] twiddle4_1_327_real;
  wire[46:0] T25040;
  wire[46:0] T25041;
  wire[46:0] T25042;
  wire[46:0] T25043;
  wire T25044;
  wire T25045;
  wire T25046;
  wire[46:0] T25047;
  wire[46:0] T25048;
  wire[46:0] T25049;
  wire[46:0] twiddle4_1_328_real;
  wire[46:0] T25050;
  wire[46:0] T25051;
  wire[46:0] T25052;
  wire[46:0] T25053;
  wire[46:0] twiddle4_1_329_real;
  wire[46:0] T25054;
  wire[46:0] T25055;
  wire[46:0] T25056;
  wire[46:0] T25057;
  wire T25058;
  wire[46:0] T25059;
  wire[46:0] twiddle4_1_330_real;
  wire[46:0] T25060;
  wire[46:0] T25061;
  wire[46:0] T25062;
  wire[46:0] T25063;
  wire[46:0] twiddle4_1_331_real;
  wire[46:0] T25064;
  wire[46:0] T25065;
  wire[46:0] T25066;
  wire[46:0] T25067;
  wire T25068;
  wire T25069;
  wire[46:0] T25070;
  wire[46:0] T25071;
  wire[46:0] twiddle4_1_332_real;
  wire[46:0] T25072;
  wire[46:0] T25073;
  wire[46:0] T25074;
  wire[46:0] T25075;
  wire[46:0] twiddle4_1_333_real;
  wire[46:0] T25076;
  wire[46:0] T25077;
  wire[46:0] T25078;
  wire[46:0] T25079;
  wire T25080;
  wire[46:0] T25081;
  wire[46:0] twiddle4_1_334_real;
  wire[46:0] T25082;
  wire[46:0] T25083;
  wire[46:0] T25084;
  wire[46:0] T25085;
  wire[46:0] twiddle4_1_335_real;
  wire[46:0] T25086;
  wire[46:0] T25087;
  wire[46:0] T25088;
  wire[46:0] T25089;
  wire T25090;
  wire T25091;
  wire T25092;
  wire T25093;
  wire[46:0] T25094;
  wire[46:0] T25095;
  wire[46:0] T25096;
  wire[46:0] T25097;
  wire[46:0] twiddle4_1_336_real;
  wire[46:0] T25098;
  wire[46:0] T25099;
  wire[46:0] T25100;
  wire[46:0] T25101;
  wire[46:0] twiddle4_1_337_real;
  wire[46:0] T25102;
  wire[46:0] T25103;
  wire[46:0] T25104;
  wire[46:0] T25105;
  wire T25106;
  wire[46:0] T25107;
  wire[46:0] twiddle4_1_338_real;
  wire[46:0] T25108;
  wire[46:0] T25109;
  wire[46:0] T25110;
  wire[46:0] T25111;
  wire[46:0] twiddle4_1_339_real;
  wire[46:0] T25112;
  wire[46:0] T25113;
  wire[46:0] T25114;
  wire[46:0] T25115;
  wire T25116;
  wire T25117;
  wire[46:0] T25118;
  wire[46:0] T25119;
  wire[46:0] twiddle4_1_340_real;
  wire[46:0] T25120;
  wire[46:0] T25121;
  wire[46:0] T25122;
  wire[46:0] T25123;
  wire[46:0] twiddle4_1_341_real;
  wire[46:0] T25124;
  wire[46:0] T25125;
  wire[46:0] T25126;
  wire[46:0] T25127;
  wire T25128;
  wire[46:0] T25129;
  wire[46:0] twiddle4_1_342_real;
  wire[46:0] T25130;
  wire[46:0] T25131;
  wire[46:0] T25132;
  wire[45:0] T25133;
  wire[45:0] T25134;
  wire T25135;
  wire[46:0] twiddle4_1_343_real;
  wire[46:0] T25136;
  wire[46:0] T25137;
  wire[46:0] T25138;
  wire[45:0] T25139;
  wire[45:0] T25140;
  wire T25141;
  wire T25142;
  wire T25143;
  wire T25144;
  wire[46:0] T25145;
  wire[46:0] T25146;
  wire[46:0] T25147;
  wire[46:0] twiddle4_1_344_real;
  wire[46:0] T25148;
  wire[46:0] T25149;
  wire[46:0] T25150;
  wire[45:0] T25151;
  wire[45:0] T25152;
  wire T25153;
  wire[46:0] twiddle4_1_345_real;
  wire[46:0] T25154;
  wire[46:0] T25155;
  wire[46:0] T25156;
  wire[45:0] T25157;
  wire[45:0] T25158;
  wire T25159;
  wire T25160;
  wire[46:0] T25161;
  wire[46:0] twiddle4_1_346_real;
  wire[46:0] T25162;
  wire[46:0] T25163;
  wire[46:0] T25164;
  wire[45:0] T25165;
  wire[45:0] T25166;
  wire T25167;
  wire[46:0] twiddle4_1_347_real;
  wire[46:0] T25168;
  wire[46:0] T25169;
  wire[46:0] T25170;
  wire[45:0] T25171;
  wire[45:0] T25172;
  wire T25173;
  wire T25174;
  wire T25175;
  wire[46:0] T25176;
  wire[46:0] T25177;
  wire[46:0] twiddle4_1_348_real;
  wire[46:0] T25178;
  wire[46:0] T25179;
  wire[46:0] T25180;
  wire[45:0] T25181;
  wire[45:0] T25182;
  wire T25183;
  wire[46:0] twiddle4_1_349_real;
  wire[46:0] T25184;
  wire[46:0] T25185;
  wire[46:0] T25186;
  wire[45:0] T25187;
  wire[45:0] T25188;
  wire T25189;
  wire T25190;
  wire[46:0] T25191;
  wire[46:0] twiddle4_1_350_real;
  wire[46:0] T25192;
  wire[46:0] T25193;
  wire[46:0] T25194;
  wire[45:0] T25195;
  wire[45:0] T25196;
  wire T25197;
  wire[46:0] twiddle4_1_351_real;
  wire[46:0] T25198;
  wire[46:0] T25199;
  wire[46:0] T25200;
  wire[45:0] T25201;
  wire[45:0] T25202;
  wire T25203;
  wire T25204;
  wire T25205;
  wire T25206;
  wire T25207;
  wire T25208;
  wire[46:0] T25209;
  wire[46:0] T25210;
  wire[46:0] T25211;
  wire[46:0] T25212;
  wire[46:0] T25213;
  wire[46:0] twiddle4_1_352_real;
  wire[46:0] T25214;
  wire[46:0] T25215;
  wire[46:0] T25216;
  wire[45:0] T25217;
  wire[45:0] T25218;
  wire T25219;
  wire[46:0] twiddle4_1_353_real;
  wire[46:0] T25220;
  wire[46:0] T25221;
  wire[46:0] T25222;
  wire[45:0] T25223;
  wire[45:0] T25224;
  wire T25225;
  wire T25226;
  wire[46:0] T25227;
  wire[46:0] twiddle4_1_354_real;
  wire[46:0] T25228;
  wire[46:0] T25229;
  wire[46:0] T25230;
  wire[45:0] T25231;
  wire[45:0] T25232;
  wire T25233;
  wire[46:0] twiddle4_1_355_real;
  wire[46:0] T25234;
  wire[46:0] T25235;
  wire[46:0] T25236;
  wire[45:0] T25237;
  wire[45:0] T25238;
  wire T25239;
  wire T25240;
  wire T25241;
  wire[46:0] T25242;
  wire[46:0] T25243;
  wire[46:0] twiddle4_1_356_real;
  wire[46:0] T25244;
  wire[46:0] T25245;
  wire[46:0] T25246;
  wire[45:0] T25247;
  wire[45:0] T25248;
  wire T25249;
  wire[46:0] twiddle4_1_357_real;
  wire[46:0] T25250;
  wire[46:0] T25251;
  wire[46:0] T25252;
  wire[45:0] T25253;
  wire[45:0] T25254;
  wire T25255;
  wire T25256;
  wire[46:0] T25257;
  wire[46:0] twiddle4_1_358_real;
  wire[46:0] T25258;
  wire[46:0] T25259;
  wire[46:0] T25260;
  wire[45:0] T25261;
  wire[45:0] T25262;
  wire T25263;
  wire[46:0] twiddle4_1_359_real;
  wire[46:0] T25264;
  wire[46:0] T25265;
  wire[46:0] T25266;
  wire[45:0] T25267;
  wire[45:0] T25268;
  wire T25269;
  wire T25270;
  wire T25271;
  wire T25272;
  wire[46:0] T25273;
  wire[46:0] T25274;
  wire[46:0] T25275;
  wire[46:0] twiddle4_1_360_real;
  wire[46:0] T25276;
  wire[46:0] T25277;
  wire[46:0] T25278;
  wire[45:0] T25279;
  wire[45:0] T25280;
  wire T25281;
  wire[46:0] twiddle4_1_361_real;
  wire[46:0] T25282;
  wire[46:0] T25283;
  wire[46:0] T25284;
  wire[45:0] T25285;
  wire[45:0] T25286;
  wire T25287;
  wire T25288;
  wire[46:0] T25289;
  wire[46:0] twiddle4_1_362_real;
  wire[46:0] T25290;
  wire[46:0] T25291;
  wire[46:0] T25292;
  wire[45:0] T25293;
  wire[45:0] T25294;
  wire T25295;
  wire[46:0] twiddle4_1_363_real;
  wire[46:0] T25296;
  wire[46:0] T25297;
  wire[46:0] T25298;
  wire[45:0] T25299;
  wire[45:0] T25300;
  wire T25301;
  wire T25302;
  wire T25303;
  wire[46:0] T25304;
  wire[46:0] T25305;
  wire[46:0] twiddle4_1_364_real;
  wire[46:0] T25306;
  wire[46:0] T25307;
  wire[46:0] T25308;
  wire[45:0] T25309;
  wire[45:0] T25310;
  wire T25311;
  wire[46:0] twiddle4_1_365_real;
  wire[46:0] T25312;
  wire[46:0] T25313;
  wire[46:0] T25314;
  wire[45:0] T25315;
  wire[45:0] T25316;
  wire T25317;
  wire T25318;
  wire[46:0] T25319;
  wire[46:0] twiddle4_1_366_real;
  wire[46:0] T25320;
  wire[46:0] T25321;
  wire[46:0] T25322;
  wire[45:0] T25323;
  wire[45:0] T25324;
  wire T25325;
  wire[46:0] twiddle4_1_367_real;
  wire[46:0] T25326;
  wire[46:0] T25327;
  wire[46:0] T25328;
  wire[45:0] T25329;
  wire[45:0] T25330;
  wire T25331;
  wire T25332;
  wire T25333;
  wire T25334;
  wire T25335;
  wire[46:0] T25336;
  wire[46:0] T25337;
  wire[46:0] T25338;
  wire[46:0] T25339;
  wire[46:0] twiddle4_1_368_real;
  wire[46:0] T25340;
  wire[46:0] T25341;
  wire[46:0] T25342;
  wire[45:0] T25343;
  wire[45:0] T25344;
  wire T25345;
  wire[46:0] twiddle4_1_369_real;
  wire[46:0] T25346;
  wire[46:0] T25347;
  wire[46:0] T25348;
  wire[45:0] T25349;
  wire[45:0] T25350;
  wire T25351;
  wire T25352;
  wire[46:0] T25353;
  wire[46:0] twiddle4_1_370_real;
  wire[46:0] T25354;
  wire[46:0] T25355;
  wire[46:0] T25356;
  wire[45:0] T25357;
  wire[45:0] T25358;
  wire T25359;
  wire[46:0] twiddle4_1_371_real;
  wire[46:0] T25360;
  wire[46:0] T25361;
  wire[46:0] T25362;
  wire[45:0] T25363;
  wire[45:0] T25364;
  wire T25365;
  wire T25366;
  wire T25367;
  wire[46:0] T25368;
  wire[46:0] T25369;
  wire[46:0] twiddle4_1_372_real;
  wire[46:0] T25370;
  wire[46:0] T25371;
  wire[46:0] T25372;
  wire[45:0] T25373;
  wire[45:0] T25374;
  wire T25375;
  wire[46:0] twiddle4_1_373_real;
  wire[46:0] T25376;
  wire[46:0] T25377;
  wire[46:0] T25378;
  wire[45:0] T25379;
  wire[45:0] T25380;
  wire T25381;
  wire T25382;
  wire[46:0] T25383;
  wire[46:0] twiddle4_1_374_real;
  wire[46:0] T25384;
  wire[46:0] T25385;
  wire[46:0] T25386;
  wire[45:0] T25387;
  wire[45:0] T25388;
  wire T25389;
  wire[46:0] twiddle4_1_375_real;
  wire[46:0] T25390;
  wire[46:0] T25391;
  wire[46:0] T25392;
  wire[45:0] T25393;
  wire[45:0] T25394;
  wire T25395;
  wire T25396;
  wire T25397;
  wire T25398;
  wire[46:0] T25399;
  wire[46:0] T25400;
  wire[46:0] T25401;
  wire[46:0] twiddle4_1_376_real;
  wire[46:0] T25402;
  wire[46:0] T25403;
  wire[46:0] T25404;
  wire[45:0] T25405;
  wire[45:0] T25406;
  wire T25407;
  wire[46:0] twiddle4_1_377_real;
  wire[46:0] T25408;
  wire[46:0] T25409;
  wire[46:0] T25410;
  wire[45:0] T25411;
  wire[45:0] T25412;
  wire T25413;
  wire T25414;
  wire[46:0] T25415;
  wire[46:0] twiddle4_1_378_real;
  wire[46:0] T25416;
  wire[46:0] T25417;
  wire[46:0] T25418;
  wire[45:0] T25419;
  wire[45:0] T25420;
  wire T25421;
  wire[46:0] twiddle4_1_379_real;
  wire[46:0] T25422;
  wire[46:0] T25423;
  wire[46:0] T25424;
  wire[45:0] T25425;
  wire[45:0] T25426;
  wire T25427;
  wire T25428;
  wire T25429;
  wire[46:0] T25430;
  wire[46:0] T25431;
  wire[46:0] twiddle4_1_380_real;
  wire[46:0] T25432;
  wire[46:0] T25433;
  wire[46:0] T25434;
  wire[45:0] T25435;
  wire[45:0] T25436;
  wire T25437;
  wire[46:0] twiddle4_1_381_real;
  wire[46:0] T25438;
  wire[46:0] T25439;
  wire[46:0] T25440;
  wire[45:0] T25441;
  wire[45:0] T25442;
  wire T25443;
  wire T25444;
  wire[46:0] T25445;
  wire[46:0] twiddle4_1_382_real;
  wire[46:0] T25446;
  wire[46:0] T25447;
  wire[46:0] T25448;
  wire[45:0] T25449;
  wire[45:0] T25450;
  wire T25451;
  wire[46:0] twiddle4_1_383_real;
  wire[46:0] T25452;
  wire[46:0] T25453;
  wire[46:0] T25454;
  wire[45:0] T25455;
  wire[45:0] T25456;
  wire T25457;
  wire T25458;
  wire T25459;
  wire T25460;
  wire T25461;
  wire T25462;
  wire T25463;
  wire T25464;
  wire[46:0] T25465;
  wire[46:0] T25466;
  wire[46:0] T25467;
  wire[46:0] T25468;
  wire[46:0] T25469;
  wire[46:0] T25470;
  wire[46:0] T25471;
  wire[46:0] twiddle4_1_384_real;
  wire[46:0] T25472;
  wire[46:0] T25473;
  wire[46:0] T25474;
  wire[45:0] T25475;
  wire[45:0] T25476;
  wire T25477;
  wire[46:0] twiddle4_1_385_real;
  wire[46:0] T25478;
  wire[46:0] T25479;
  wire[46:0] T25480;
  wire[45:0] T25481;
  wire[45:0] T25482;
  wire T25483;
  wire T25484;
  wire[46:0] T25485;
  wire[46:0] twiddle4_1_386_real;
  wire[46:0] T25486;
  wire[46:0] T25487;
  wire[46:0] T25488;
  wire[45:0] T25489;
  wire[45:0] T25490;
  wire T25491;
  wire[46:0] twiddle4_1_387_real;
  wire[46:0] T25492;
  wire[46:0] T25493;
  wire[46:0] T25494;
  wire[45:0] T25495;
  wire[45:0] T25496;
  wire T25497;
  wire T25498;
  wire T25499;
  wire[46:0] T25500;
  wire[46:0] T25501;
  wire[46:0] twiddle4_1_388_real;
  wire[46:0] T25502;
  wire[46:0] T25503;
  wire[46:0] T25504;
  wire[45:0] T25505;
  wire[45:0] T25506;
  wire T25507;
  wire[46:0] twiddle4_1_389_real;
  wire[46:0] T25508;
  wire[46:0] T25509;
  wire[46:0] T25510;
  wire[45:0] T25511;
  wire[45:0] T25512;
  wire T25513;
  wire T25514;
  wire[46:0] T25515;
  wire[46:0] twiddle4_1_390_real;
  wire[46:0] T25516;
  wire[46:0] T25517;
  wire[46:0] T25518;
  wire[45:0] T25519;
  wire[45:0] T25520;
  wire T25521;
  wire[46:0] twiddle4_1_391_real;
  wire[46:0] T25522;
  wire[46:0] T25523;
  wire[46:0] T25524;
  wire[45:0] T25525;
  wire[45:0] T25526;
  wire T25527;
  wire T25528;
  wire T25529;
  wire T25530;
  wire[46:0] T25531;
  wire[46:0] T25532;
  wire[46:0] T25533;
  wire[46:0] twiddle4_1_392_real;
  wire[46:0] T25534;
  wire[46:0] T25535;
  wire[46:0] T25536;
  wire[45:0] T25537;
  wire[45:0] T25538;
  wire T25539;
  wire[46:0] twiddle4_1_393_real;
  wire[46:0] T25540;
  wire[46:0] T25541;
  wire[46:0] T25542;
  wire[45:0] T25543;
  wire[45:0] T25544;
  wire T25545;
  wire T25546;
  wire[46:0] T25547;
  wire[46:0] twiddle4_1_394_real;
  wire[46:0] T25548;
  wire[46:0] T25549;
  wire[46:0] T25550;
  wire[45:0] T25551;
  wire[45:0] T25552;
  wire T25553;
  wire[46:0] twiddle4_1_395_real;
  wire[46:0] T25554;
  wire[46:0] T25555;
  wire[46:0] T25556;
  wire[45:0] T25557;
  wire[45:0] T25558;
  wire T25559;
  wire T25560;
  wire T25561;
  wire[46:0] T25562;
  wire[46:0] T25563;
  wire[46:0] twiddle4_1_396_real;
  wire[46:0] T25564;
  wire[46:0] T25565;
  wire[46:0] T25566;
  wire[45:0] T25567;
  wire[45:0] T25568;
  wire T25569;
  wire[46:0] twiddle4_1_397_real;
  wire[46:0] T25570;
  wire[46:0] T25571;
  wire[46:0] T25572;
  wire[45:0] T25573;
  wire[45:0] T25574;
  wire T25575;
  wire T25576;
  wire[46:0] T25577;
  wire[46:0] twiddle4_1_398_real;
  wire[46:0] T25578;
  wire[46:0] T25579;
  wire[46:0] T25580;
  wire[45:0] T25581;
  wire[45:0] T25582;
  wire T25583;
  wire[46:0] twiddle4_1_399_real;
  wire[46:0] T25584;
  wire[46:0] T25585;
  wire[46:0] T25586;
  wire[45:0] T25587;
  wire[45:0] T25588;
  wire T25589;
  wire T25590;
  wire T25591;
  wire T25592;
  wire T25593;
  wire[46:0] T25594;
  wire[46:0] T25595;
  wire[46:0] T25596;
  wire[46:0] T25597;
  wire[46:0] twiddle4_1_400_real;
  wire[46:0] T25598;
  wire[46:0] T25599;
  wire[46:0] T25600;
  wire[45:0] T25601;
  wire[45:0] T25602;
  wire T25603;
  wire[46:0] twiddle4_1_401_real;
  wire[46:0] T25604;
  wire[46:0] T25605;
  wire[46:0] T25606;
  wire[45:0] T25607;
  wire[45:0] T25608;
  wire T25609;
  wire T25610;
  wire[46:0] T25611;
  wire[46:0] twiddle4_1_402_real;
  wire[46:0] T25612;
  wire[46:0] T25613;
  wire[46:0] T25614;
  wire[45:0] T25615;
  wire[45:0] T25616;
  wire T25617;
  wire[46:0] twiddle4_1_403_real;
  wire[46:0] T25618;
  wire[46:0] T25619;
  wire[46:0] T25620;
  wire[45:0] T25621;
  wire[45:0] T25622;
  wire T25623;
  wire T25624;
  wire T25625;
  wire[46:0] T25626;
  wire[46:0] T25627;
  wire[46:0] twiddle4_1_404_real;
  wire[46:0] T25628;
  wire[46:0] T25629;
  wire[46:0] T25630;
  wire[45:0] T25631;
  wire[45:0] T25632;
  wire T25633;
  wire[46:0] twiddle4_1_405_real;
  wire[46:0] T25634;
  wire[46:0] T25635;
  wire[46:0] T25636;
  wire[45:0] T25637;
  wire[45:0] T25638;
  wire T25639;
  wire T25640;
  wire[46:0] T25641;
  wire[46:0] twiddle4_1_406_real;
  wire[46:0] T25642;
  wire[46:0] T25643;
  wire[46:0] T25644;
  wire[45:0] T25645;
  wire[45:0] T25646;
  wire T25647;
  wire[46:0] twiddle4_1_407_real;
  wire[46:0] T25648;
  wire[46:0] T25649;
  wire[46:0] T25650;
  wire[45:0] T25651;
  wire[45:0] T25652;
  wire T25653;
  wire T25654;
  wire T25655;
  wire T25656;
  wire[46:0] T25657;
  wire[46:0] T25658;
  wire[46:0] T25659;
  wire[46:0] twiddle4_1_408_real;
  wire[46:0] T25660;
  wire[46:0] T25661;
  wire[46:0] T25662;
  wire[45:0] T25663;
  wire[45:0] T25664;
  wire T25665;
  wire[46:0] twiddle4_1_409_real;
  wire[46:0] T25666;
  wire[46:0] T25667;
  wire[46:0] T25668;
  wire[45:0] T25669;
  wire[45:0] T25670;
  wire T25671;
  wire T25672;
  wire[46:0] T25673;
  wire[46:0] twiddle4_1_410_real;
  wire[46:0] T25674;
  wire[46:0] T25675;
  wire[46:0] T25676;
  wire[45:0] T25677;
  wire[45:0] T25678;
  wire T25679;
  wire[46:0] twiddle4_1_411_real;
  wire[46:0] T25680;
  wire[46:0] T25681;
  wire[46:0] T25682;
  wire[45:0] T25683;
  wire[45:0] T25684;
  wire T25685;
  wire T25686;
  wire T25687;
  wire[46:0] T25688;
  wire[46:0] T25689;
  wire[46:0] twiddle4_1_412_real;
  wire[46:0] T25690;
  wire[46:0] T25691;
  wire[46:0] T25692;
  wire[45:0] T25693;
  wire[45:0] T25694;
  wire T25695;
  wire[46:0] twiddle4_1_413_real;
  wire[46:0] T25696;
  wire[46:0] T25697;
  wire[46:0] T25698;
  wire[45:0] T25699;
  wire[45:0] T25700;
  wire T25701;
  wire T25702;
  wire[46:0] T25703;
  wire[46:0] twiddle4_1_414_real;
  wire[46:0] T25704;
  wire[46:0] T25705;
  wire[46:0] T25706;
  wire[45:0] T25707;
  wire[45:0] T25708;
  wire T25709;
  wire[46:0] twiddle4_1_415_real;
  wire[46:0] T25710;
  wire[46:0] T25711;
  wire[46:0] T25712;
  wire[45:0] T25713;
  wire[45:0] T25714;
  wire T25715;
  wire T25716;
  wire T25717;
  wire T25718;
  wire T25719;
  wire T25720;
  wire[46:0] T25721;
  wire[46:0] T25722;
  wire[46:0] T25723;
  wire[46:0] T25724;
  wire[46:0] T25725;
  wire[46:0] twiddle4_1_416_real;
  wire[46:0] T25726;
  wire[46:0] T25727;
  wire[46:0] T25728;
  wire[45:0] T25729;
  wire[45:0] T25730;
  wire T25731;
  wire[46:0] twiddle4_1_417_real;
  wire[46:0] T25732;
  wire[46:0] T25733;
  wire[46:0] T25734;
  wire[45:0] T25735;
  wire[45:0] T25736;
  wire T25737;
  wire T25738;
  wire[46:0] T25739;
  wire[46:0] twiddle4_1_418_real;
  wire[46:0] T25740;
  wire[46:0] T25741;
  wire[46:0] T25742;
  wire[45:0] T25743;
  wire[45:0] T25744;
  wire T25745;
  wire[46:0] twiddle4_1_419_real;
  wire[46:0] T25746;
  wire[46:0] T25747;
  wire[46:0] T25748;
  wire[45:0] T25749;
  wire[45:0] T25750;
  wire T25751;
  wire T25752;
  wire T25753;
  wire[46:0] T25754;
  wire[46:0] T25755;
  wire[46:0] twiddle4_1_420_real;
  wire[46:0] T25756;
  wire[46:0] T25757;
  wire[46:0] T25758;
  wire[45:0] T25759;
  wire[45:0] T25760;
  wire T25761;
  wire[46:0] twiddle4_1_421_real;
  wire[46:0] T25762;
  wire[46:0] T25763;
  wire[46:0] T25764;
  wire[45:0] T25765;
  wire[45:0] T25766;
  wire T25767;
  wire T25768;
  wire[46:0] T25769;
  wire[46:0] twiddle4_1_422_real;
  wire[46:0] T25770;
  wire[46:0] T25771;
  wire[46:0] T25772;
  wire[45:0] T25773;
  wire[45:0] T25774;
  wire T25775;
  wire[46:0] twiddle4_1_423_real;
  wire[46:0] T25776;
  wire[46:0] T25777;
  wire[46:0] T25778;
  wire[45:0] T25779;
  wire[45:0] T25780;
  wire T25781;
  wire T25782;
  wire T25783;
  wire T25784;
  wire[46:0] T25785;
  wire[46:0] T25786;
  wire[46:0] T25787;
  wire[46:0] twiddle4_1_424_real;
  wire[46:0] T25788;
  wire[46:0] T25789;
  wire[46:0] T25790;
  wire[45:0] T25791;
  wire[45:0] T25792;
  wire T25793;
  wire[46:0] twiddle4_1_425_real;
  wire[46:0] T25794;
  wire[46:0] T25795;
  wire[46:0] T25796;
  wire[45:0] T25797;
  wire[45:0] T25798;
  wire T25799;
  wire T25800;
  wire[46:0] T25801;
  wire[46:0] twiddle4_1_426_real;
  wire[46:0] T25802;
  wire[46:0] T25803;
  wire[46:0] T25804;
  wire[45:0] T25805;
  wire[45:0] T25806;
  wire T25807;
  wire[46:0] twiddle4_1_427_real;
  wire[46:0] T25808;
  wire[46:0] T25809;
  wire[46:0] T25810;
  wire[45:0] T25811;
  wire[45:0] T25812;
  wire T25813;
  wire T25814;
  wire T25815;
  wire[46:0] T25816;
  wire[46:0] T25817;
  wire[46:0] twiddle4_1_428_real;
  wire[46:0] T25818;
  wire[46:0] T25819;
  wire[46:0] T25820;
  wire[45:0] T25821;
  wire[45:0] T25822;
  wire T25823;
  wire[46:0] twiddle4_1_429_real;
  wire[46:0] T25824;
  wire[46:0] T25825;
  wire[46:0] T25826;
  wire[45:0] T25827;
  wire[45:0] T25828;
  wire T25829;
  wire T25830;
  wire[46:0] T25831;
  wire[46:0] twiddle4_1_430_real;
  wire[46:0] T25832;
  wire[46:0] T25833;
  wire[46:0] T25834;
  wire[44:0] T25835;
  wire[44:0] T25836;
  wire[1:0] T25837;
  wire T25838;
  wire[46:0] twiddle4_1_431_real;
  wire[46:0] T25839;
  wire[46:0] T25840;
  wire[46:0] T25841;
  wire[44:0] T25842;
  wire[44:0] T25843;
  wire[1:0] T25844;
  wire T25845;
  wire T25846;
  wire T25847;
  wire T25848;
  wire T25849;
  wire[46:0] T25850;
  wire[46:0] T25851;
  wire[46:0] T25852;
  wire[46:0] T25853;
  wire[46:0] twiddle4_1_432_real;
  wire[46:0] T25854;
  wire[46:0] T25855;
  wire[46:0] T25856;
  wire[44:0] T25857;
  wire[44:0] T25858;
  wire[1:0] T25859;
  wire T25860;
  wire[46:0] twiddle4_1_433_real;
  wire[46:0] T25861;
  wire[46:0] T25862;
  wire[46:0] T25863;
  wire[44:0] T25864;
  wire[44:0] T25865;
  wire[1:0] T25866;
  wire T25867;
  wire T25868;
  wire[46:0] T25869;
  wire[46:0] twiddle4_1_434_real;
  wire[46:0] T25870;
  wire[46:0] T25871;
  wire[46:0] T25872;
  wire[44:0] T25873;
  wire[44:0] T25874;
  wire[1:0] T25875;
  wire T25876;
  wire[46:0] twiddle4_1_435_real;
  wire[46:0] T25877;
  wire[46:0] T25878;
  wire[46:0] T25879;
  wire[44:0] T25880;
  wire[44:0] T25881;
  wire[1:0] T25882;
  wire T25883;
  wire T25884;
  wire T25885;
  wire[46:0] T25886;
  wire[46:0] T25887;
  wire[46:0] twiddle4_1_436_real;
  wire[46:0] T25888;
  wire[46:0] T25889;
  wire[46:0] T25890;
  wire[44:0] T25891;
  wire[44:0] T25892;
  wire[1:0] T25893;
  wire T25894;
  wire[46:0] twiddle4_1_437_real;
  wire[46:0] T25895;
  wire[46:0] T25896;
  wire[46:0] T25897;
  wire[44:0] T25898;
  wire[44:0] T25899;
  wire[1:0] T25900;
  wire T25901;
  wire T25902;
  wire[46:0] T25903;
  wire[46:0] twiddle4_1_438_real;
  wire[46:0] T25904;
  wire[46:0] T25905;
  wire[46:0] T25906;
  wire[44:0] T25907;
  wire[44:0] T25908;
  wire[1:0] T25909;
  wire T25910;
  wire[46:0] twiddle4_1_439_real;
  wire[46:0] T25911;
  wire[46:0] T25912;
  wire[46:0] T25913;
  wire[44:0] T25914;
  wire[44:0] T25915;
  wire[1:0] T25916;
  wire T25917;
  wire T25918;
  wire T25919;
  wire T25920;
  wire[46:0] T25921;
  wire[46:0] T25922;
  wire[46:0] T25923;
  wire[46:0] twiddle4_1_440_real;
  wire[46:0] T25924;
  wire[46:0] T25925;
  wire[46:0] T25926;
  wire[44:0] T25927;
  wire[44:0] T25928;
  wire[1:0] T25929;
  wire T25930;
  wire[46:0] twiddle4_1_441_real;
  wire[46:0] T25931;
  wire[46:0] T25932;
  wire[46:0] T25933;
  wire[44:0] T25934;
  wire[44:0] T25935;
  wire[1:0] T25936;
  wire T25937;
  wire T25938;
  wire[46:0] T25939;
  wire[46:0] twiddle4_1_442_real;
  wire[46:0] T25940;
  wire[46:0] T25941;
  wire[46:0] T25942;
  wire[44:0] T25943;
  wire[44:0] T25944;
  wire[1:0] T25945;
  wire T25946;
  wire[46:0] twiddle4_1_443_real;
  wire[46:0] T25947;
  wire[46:0] T25948;
  wire[46:0] T25949;
  wire[44:0] T25950;
  wire[44:0] T25951;
  wire[1:0] T25952;
  wire T25953;
  wire T25954;
  wire T25955;
  wire[46:0] T25956;
  wire[46:0] T25957;
  wire[46:0] twiddle4_1_444_real;
  wire[46:0] T25958;
  wire[46:0] T25959;
  wire[46:0] T25960;
  wire[44:0] T25961;
  wire[44:0] T25962;
  wire[1:0] T25963;
  wire T25964;
  wire[46:0] twiddle4_1_445_real;
  wire[46:0] T25965;
  wire[46:0] T25966;
  wire[46:0] T25967;
  wire[44:0] T25968;
  wire[44:0] T25969;
  wire[1:0] T25970;
  wire T25971;
  wire T25972;
  wire[46:0] T25973;
  wire[46:0] twiddle4_1_446_real;
  wire[46:0] T25974;
  wire[46:0] T25975;
  wire[46:0] T25976;
  wire[44:0] T25977;
  wire[44:0] T25978;
  wire[1:0] T25979;
  wire T25980;
  wire[46:0] twiddle4_1_447_real;
  wire[46:0] T25981;
  wire[46:0] T25982;
  wire[46:0] T25983;
  wire[44:0] T25984;
  wire[44:0] T25985;
  wire[1:0] T25986;
  wire T25987;
  wire T25988;
  wire T25989;
  wire T25990;
  wire T25991;
  wire T25992;
  wire T25993;
  wire[46:0] T25994;
  wire[46:0] T25995;
  wire[46:0] T25996;
  wire[46:0] T25997;
  wire[46:0] T25998;
  wire[46:0] T25999;
  wire[46:0] twiddle4_1_448_real;
  wire[46:0] T26000;
  wire[46:0] T26001;
  wire[46:0] T26002;
  wire[44:0] T26003;
  wire[44:0] T26004;
  wire[1:0] T26005;
  wire T26006;
  wire[46:0] twiddle4_1_449_real;
  wire[46:0] T26007;
  wire[46:0] T26008;
  wire[46:0] T26009;
  wire[44:0] T26010;
  wire[44:0] T26011;
  wire[1:0] T26012;
  wire T26013;
  wire T26014;
  wire[46:0] T26015;
  wire[46:0] twiddle4_1_450_real;
  wire[46:0] T26016;
  wire[46:0] T26017;
  wire[46:0] T26018;
  wire[44:0] T26019;
  wire[44:0] T26020;
  wire[1:0] T26021;
  wire T26022;
  wire[46:0] twiddle4_1_451_real;
  wire[46:0] T26023;
  wire[46:0] T26024;
  wire[46:0] T26025;
  wire[44:0] T26026;
  wire[44:0] T26027;
  wire[1:0] T26028;
  wire T26029;
  wire T26030;
  wire T26031;
  wire[46:0] T26032;
  wire[46:0] T26033;
  wire[46:0] twiddle4_1_452_real;
  wire[46:0] T26034;
  wire[46:0] T26035;
  wire[46:0] T26036;
  wire[44:0] T26037;
  wire[44:0] T26038;
  wire[1:0] T26039;
  wire T26040;
  wire[46:0] twiddle4_1_453_real;
  wire[46:0] T26041;
  wire[46:0] T26042;
  wire[46:0] T26043;
  wire[44:0] T26044;
  wire[44:0] T26045;
  wire[1:0] T26046;
  wire T26047;
  wire T26048;
  wire[46:0] T26049;
  wire[46:0] twiddle4_1_454_real;
  wire[46:0] T26050;
  wire[46:0] T26051;
  wire[46:0] T26052;
  wire[44:0] T26053;
  wire[44:0] T26054;
  wire[1:0] T26055;
  wire T26056;
  wire[46:0] twiddle4_1_455_real;
  wire[46:0] T26057;
  wire[46:0] T26058;
  wire[46:0] T26059;
  wire[44:0] T26060;
  wire[44:0] T26061;
  wire[1:0] T26062;
  wire T26063;
  wire T26064;
  wire T26065;
  wire T26066;
  wire[46:0] T26067;
  wire[46:0] T26068;
  wire[46:0] T26069;
  wire[46:0] twiddle4_1_456_real;
  wire[46:0] T26070;
  wire[46:0] T26071;
  wire[46:0] T26072;
  wire[44:0] T26073;
  wire[44:0] T26074;
  wire[1:0] T26075;
  wire T26076;
  wire[46:0] twiddle4_1_457_real;
  wire[46:0] T26077;
  wire[46:0] T26078;
  wire[46:0] T26079;
  wire[44:0] T26080;
  wire[44:0] T26081;
  wire[1:0] T26082;
  wire T26083;
  wire T26084;
  wire[46:0] T26085;
  wire[46:0] twiddle4_1_458_real;
  wire[46:0] T26086;
  wire[46:0] T26087;
  wire[46:0] T26088;
  wire[44:0] T26089;
  wire[44:0] T26090;
  wire[1:0] T26091;
  wire T26092;
  wire[46:0] twiddle4_1_459_real;
  wire[46:0] T26093;
  wire[46:0] T26094;
  wire[46:0] T26095;
  wire[44:0] T26096;
  wire[44:0] T26097;
  wire[1:0] T26098;
  wire T26099;
  wire T26100;
  wire T26101;
  wire[46:0] T26102;
  wire[46:0] T26103;
  wire[46:0] twiddle4_1_460_real;
  wire[46:0] T26104;
  wire[46:0] T26105;
  wire[46:0] T26106;
  wire[44:0] T26107;
  wire[44:0] T26108;
  wire[1:0] T26109;
  wire T26110;
  wire[46:0] twiddle4_1_461_real;
  wire[46:0] T26111;
  wire[46:0] T26112;
  wire[46:0] T26113;
  wire[44:0] T26114;
  wire[44:0] T26115;
  wire[1:0] T26116;
  wire T26117;
  wire T26118;
  wire[46:0] T26119;
  wire[46:0] twiddle4_1_462_real;
  wire[46:0] T26120;
  wire[46:0] T26121;
  wire[46:0] T26122;
  wire[44:0] T26123;
  wire[44:0] T26124;
  wire[1:0] T26125;
  wire T26126;
  wire[46:0] twiddle4_1_463_real;
  wire[46:0] T26127;
  wire[46:0] T26128;
  wire[46:0] T26129;
  wire[44:0] T26130;
  wire[44:0] T26131;
  wire[1:0] T26132;
  wire T26133;
  wire T26134;
  wire T26135;
  wire T26136;
  wire T26137;
  wire[46:0] T26138;
  wire[46:0] T26139;
  wire[46:0] T26140;
  wire[46:0] T26141;
  wire[46:0] twiddle4_1_464_real;
  wire[46:0] T26142;
  wire[46:0] T26143;
  wire[46:0] T26144;
  wire[44:0] T26145;
  wire[44:0] T26146;
  wire[1:0] T26147;
  wire T26148;
  wire[46:0] twiddle4_1_465_real;
  wire[46:0] T26149;
  wire[46:0] T26150;
  wire[46:0] T26151;
  wire[44:0] T26152;
  wire[44:0] T26153;
  wire[1:0] T26154;
  wire T26155;
  wire T26156;
  wire[46:0] T26157;
  wire[46:0] twiddle4_1_466_real;
  wire[46:0] T26158;
  wire[46:0] T26159;
  wire[46:0] T26160;
  wire[44:0] T26161;
  wire[44:0] T26162;
  wire[1:0] T26163;
  wire T26164;
  wire[46:0] twiddle4_1_467_real;
  wire[46:0] T26165;
  wire[46:0] T26166;
  wire[46:0] T26167;
  wire[44:0] T26168;
  wire[44:0] T26169;
  wire[1:0] T26170;
  wire T26171;
  wire T26172;
  wire T26173;
  wire[46:0] T26174;
  wire[46:0] T26175;
  wire[46:0] twiddle4_1_468_real;
  wire[46:0] T26176;
  wire[46:0] T26177;
  wire[46:0] T26178;
  wire[44:0] T26179;
  wire[44:0] T26180;
  wire[1:0] T26181;
  wire T26182;
  wire[46:0] twiddle4_1_469_real;
  wire[46:0] T26183;
  wire[46:0] T26184;
  wire[46:0] T26185;
  wire[44:0] T26186;
  wire[44:0] T26187;
  wire[1:0] T26188;
  wire T26189;
  wire T26190;
  wire[46:0] T26191;
  wire[46:0] twiddle4_1_470_real;
  wire[46:0] T26192;
  wire[46:0] T26193;
  wire[46:0] T26194;
  wire[44:0] T26195;
  wire[44:0] T26196;
  wire[1:0] T26197;
  wire T26198;
  wire[46:0] twiddle4_1_471_real;
  wire[46:0] T26199;
  wire[46:0] T26200;
  wire[46:0] T26201;
  wire[44:0] T26202;
  wire[44:0] T26203;
  wire[1:0] T26204;
  wire T26205;
  wire T26206;
  wire T26207;
  wire T26208;
  wire[46:0] T26209;
  wire[46:0] T26210;
  wire[46:0] T26211;
  wire[46:0] twiddle4_1_472_real;
  wire[46:0] T26212;
  wire[46:0] T26213;
  wire[46:0] T26214;
  wire[43:0] T26215;
  wire[43:0] T26216;
  wire[2:0] T26217;
  wire T26218;
  wire[46:0] twiddle4_1_473_real;
  wire[46:0] T26219;
  wire[46:0] T26220;
  wire[46:0] T26221;
  wire[43:0] T26222;
  wire[43:0] T26223;
  wire[2:0] T26224;
  wire T26225;
  wire T26226;
  wire[46:0] T26227;
  wire[46:0] twiddle4_1_474_real;
  wire[46:0] T26228;
  wire[46:0] T26229;
  wire[46:0] T26230;
  wire[43:0] T26231;
  wire[43:0] T26232;
  wire[2:0] T26233;
  wire T26234;
  wire[46:0] twiddle4_1_475_real;
  wire[46:0] T26235;
  wire[46:0] T26236;
  wire[46:0] T26237;
  wire[43:0] T26238;
  wire[43:0] T26239;
  wire[2:0] T26240;
  wire T26241;
  wire T26242;
  wire T26243;
  wire[46:0] T26244;
  wire[46:0] T26245;
  wire[46:0] twiddle4_1_476_real;
  wire[46:0] T26246;
  wire[46:0] T26247;
  wire[46:0] T26248;
  wire[43:0] T26249;
  wire[43:0] T26250;
  wire[2:0] T26251;
  wire T26252;
  wire[46:0] twiddle4_1_477_real;
  wire[46:0] T26253;
  wire[46:0] T26254;
  wire[46:0] T26255;
  wire[43:0] T26256;
  wire[43:0] T26257;
  wire[2:0] T26258;
  wire T26259;
  wire T26260;
  wire[46:0] T26261;
  wire[46:0] twiddle4_1_478_real;
  wire[46:0] T26262;
  wire[46:0] T26263;
  wire[46:0] T26264;
  wire[43:0] T26265;
  wire[43:0] T26266;
  wire[2:0] T26267;
  wire T26268;
  wire[46:0] twiddle4_1_479_real;
  wire[46:0] T26269;
  wire[46:0] T26270;
  wire[46:0] T26271;
  wire[43:0] T26272;
  wire[43:0] T26273;
  wire[2:0] T26274;
  wire T26275;
  wire T26276;
  wire T26277;
  wire T26278;
  wire T26279;
  wire T26280;
  wire[46:0] T26281;
  wire[46:0] T26282;
  wire[46:0] T26283;
  wire[46:0] T26284;
  wire[46:0] T26285;
  wire[46:0] twiddle4_1_480_real;
  wire[46:0] T26286;
  wire[46:0] T26287;
  wire[46:0] T26288;
  wire[43:0] T26289;
  wire[43:0] T26290;
  wire[2:0] T26291;
  wire T26292;
  wire[46:0] twiddle4_1_481_real;
  wire[46:0] T26293;
  wire[46:0] T26294;
  wire[46:0] T26295;
  wire[43:0] T26296;
  wire[43:0] T26297;
  wire[2:0] T26298;
  wire T26299;
  wire T26300;
  wire[46:0] T26301;
  wire[46:0] twiddle4_1_482_real;
  wire[46:0] T26302;
  wire[46:0] T26303;
  wire[46:0] T26304;
  wire[43:0] T26305;
  wire[43:0] T26306;
  wire[2:0] T26307;
  wire T26308;
  wire[46:0] twiddle4_1_483_real;
  wire[46:0] T26309;
  wire[46:0] T26310;
  wire[46:0] T26311;
  wire[43:0] T26312;
  wire[43:0] T26313;
  wire[2:0] T26314;
  wire T26315;
  wire T26316;
  wire T26317;
  wire[46:0] T26318;
  wire[46:0] T26319;
  wire[46:0] twiddle4_1_484_real;
  wire[46:0] T26320;
  wire[46:0] T26321;
  wire[46:0] T26322;
  wire[43:0] T26323;
  wire[43:0] T26324;
  wire[2:0] T26325;
  wire T26326;
  wire[46:0] twiddle4_1_485_real;
  wire[46:0] T26327;
  wire[46:0] T26328;
  wire[46:0] T26329;
  wire[43:0] T26330;
  wire[43:0] T26331;
  wire[2:0] T26332;
  wire T26333;
  wire T26334;
  wire[46:0] T26335;
  wire[46:0] twiddle4_1_486_real;
  wire[46:0] T26336;
  wire[46:0] T26337;
  wire[46:0] T26338;
  wire[43:0] T26339;
  wire[43:0] T26340;
  wire[2:0] T26341;
  wire T26342;
  wire[46:0] twiddle4_1_487_real;
  wire[46:0] T26343;
  wire[46:0] T26344;
  wire[46:0] T26345;
  wire[43:0] T26346;
  wire[43:0] T26347;
  wire[2:0] T26348;
  wire T26349;
  wire T26350;
  wire T26351;
  wire T26352;
  wire[46:0] T26353;
  wire[46:0] T26354;
  wire[46:0] T26355;
  wire[46:0] twiddle4_1_488_real;
  wire[46:0] T26356;
  wire[46:0] T26357;
  wire[46:0] T26358;
  wire[43:0] T26359;
  wire[43:0] T26360;
  wire[2:0] T26361;
  wire T26362;
  wire[46:0] twiddle4_1_489_real;
  wire[46:0] T26363;
  wire[46:0] T26364;
  wire[46:0] T26365;
  wire[43:0] T26366;
  wire[43:0] T26367;
  wire[2:0] T26368;
  wire T26369;
  wire T26370;
  wire[46:0] T26371;
  wire[46:0] twiddle4_1_490_real;
  wire[46:0] T26372;
  wire[46:0] T26373;
  wire[46:0] T26374;
  wire[43:0] T26375;
  wire[43:0] T26376;
  wire[2:0] T26377;
  wire T26378;
  wire[46:0] twiddle4_1_491_real;
  wire[46:0] T26379;
  wire[46:0] T26380;
  wire[46:0] T26381;
  wire[43:0] T26382;
  wire[43:0] T26383;
  wire[2:0] T26384;
  wire T26385;
  wire T26386;
  wire T26387;
  wire[46:0] T26388;
  wire[46:0] T26389;
  wire[46:0] twiddle4_1_492_real;
  wire[46:0] T26390;
  wire[46:0] T26391;
  wire[46:0] T26392;
  wire[42:0] T26393;
  wire[42:0] T26394;
  wire[3:0] T26395;
  wire T26396;
  wire[46:0] twiddle4_1_493_real;
  wire[46:0] T26397;
  wire[46:0] T26398;
  wire[46:0] T26399;
  wire[42:0] T26400;
  wire[42:0] T26401;
  wire[3:0] T26402;
  wire T26403;
  wire T26404;
  wire[46:0] T26405;
  wire[46:0] twiddle4_1_494_real;
  wire[46:0] T26406;
  wire[46:0] T26407;
  wire[46:0] T26408;
  wire[42:0] T26409;
  wire[42:0] T26410;
  wire[3:0] T26411;
  wire T26412;
  wire[46:0] twiddle4_1_495_real;
  wire[46:0] T26413;
  wire[46:0] T26414;
  wire[46:0] T26415;
  wire[42:0] T26416;
  wire[42:0] T26417;
  wire[3:0] T26418;
  wire T26419;
  wire T26420;
  wire T26421;
  wire T26422;
  wire T26423;
  wire[46:0] T26424;
  wire[46:0] T26425;
  wire[46:0] T26426;
  wire[46:0] T26427;
  wire[46:0] twiddle4_1_496_real;
  wire[46:0] T26428;
  wire[46:0] T26429;
  wire[46:0] T26430;
  wire[42:0] T26431;
  wire[42:0] T26432;
  wire[3:0] T26433;
  wire T26434;
  wire[46:0] twiddle4_1_497_real;
  wire[46:0] T26435;
  wire[46:0] T26436;
  wire[46:0] T26437;
  wire[42:0] T26438;
  wire[42:0] T26439;
  wire[3:0] T26440;
  wire T26441;
  wire T26442;
  wire[46:0] T26443;
  wire[46:0] twiddle4_1_498_real;
  wire[46:0] T26444;
  wire[46:0] T26445;
  wire[46:0] T26446;
  wire[42:0] T26447;
  wire[42:0] T26448;
  wire[3:0] T26449;
  wire T26450;
  wire[46:0] twiddle4_1_499_real;
  wire[46:0] T26451;
  wire[46:0] T26452;
  wire[46:0] T26453;
  wire[42:0] T26454;
  wire[42:0] T26455;
  wire[3:0] T26456;
  wire T26457;
  wire T26458;
  wire T26459;
  wire[46:0] T26460;
  wire[46:0] T26461;
  wire[46:0] twiddle4_1_500_real;
  wire[46:0] T26462;
  wire[46:0] T26463;
  wire[46:0] T26464;
  wire[42:0] T26465;
  wire[42:0] T26466;
  wire[3:0] T26467;
  wire T26468;
  wire[46:0] twiddle4_1_501_real;
  wire[46:0] T26469;
  wire[46:0] T26470;
  wire[46:0] T26471;
  wire[42:0] T26472;
  wire[42:0] T26473;
  wire[3:0] T26474;
  wire T26475;
  wire T26476;
  wire[46:0] T26477;
  wire[46:0] twiddle4_1_502_real;
  wire[46:0] T26478;
  wire[46:0] T26479;
  wire[46:0] T26480;
  wire[41:0] T26481;
  wire[41:0] T26482;
  wire[4:0] T26483;
  wire T26484;
  wire[46:0] twiddle4_1_503_real;
  wire[46:0] T26485;
  wire[46:0] T26486;
  wire[46:0] T26487;
  wire[41:0] T26488;
  wire[41:0] T26489;
  wire[4:0] T26490;
  wire T26491;
  wire T26492;
  wire T26493;
  wire T26494;
  wire[46:0] T26495;
  wire[46:0] T26496;
  wire[46:0] T26497;
  wire[46:0] twiddle4_1_504_real;
  wire[46:0] T26498;
  wire[46:0] T26499;
  wire[46:0] T26500;
  wire[41:0] T26501;
  wire[41:0] T26502;
  wire[4:0] T26503;
  wire T26504;
  wire[46:0] twiddle4_1_505_real;
  wire[46:0] T26505;
  wire[46:0] T26506;
  wire[46:0] T26507;
  wire[41:0] T26508;
  wire[41:0] T26509;
  wire[4:0] T26510;
  wire T26511;
  wire T26512;
  wire[46:0] T26513;
  wire[46:0] twiddle4_1_506_real;
  wire[46:0] T26514;
  wire[46:0] T26515;
  wire[46:0] T26516;
  wire[41:0] T26517;
  wire[41:0] T26518;
  wire[4:0] T26519;
  wire T26520;
  wire[46:0] twiddle4_1_507_real;
  wire[46:0] T26521;
  wire[46:0] T26522;
  wire[46:0] T26523;
  wire[40:0] T26524;
  wire[40:0] T26525;
  wire[5:0] T26526;
  wire T26527;
  wire T26528;
  wire T26529;
  wire[46:0] T26530;
  wire[46:0] T26531;
  wire[46:0] twiddle4_1_508_real;
  wire[46:0] T26532;
  wire[46:0] T26533;
  wire[46:0] T26534;
  wire[40:0] T26535;
  wire[40:0] T26536;
  wire[5:0] T26537;
  wire T26538;
  wire[46:0] twiddle4_1_509_real;
  wire[46:0] T26539;
  wire[46:0] T26540;
  wire[46:0] T26541;
  wire[40:0] T26542;
  wire[40:0] T26543;
  wire[5:0] T26544;
  wire T26545;
  wire T26546;
  wire[46:0] T26547;
  wire[46:0] twiddle4_1_510_real;
  wire[46:0] T26548;
  wire[46:0] T26549;
  wire[46:0] T26550;
  wire[39:0] T26551;
  wire[39:0] T26552;
  wire[6:0] T26553;
  wire T26554;
  wire[46:0] twiddle4_1_511_real;
  wire[46:0] T26555;
  wire[46:0] T26556;
  wire[46:0] T26557;
  wire[38:0] T26558;
  wire[38:0] T26559;
  wire[7:0] T26560;
  wire T26561;
  wire T26562;
  wire T26563;
  wire T26564;
  wire T26565;
  wire T26566;
  wire T26567;
  wire T26568;
  wire T26569;
  wire T26570;
  wire T26571;


  assign io_t5_4out_imag = T0;
  assign T0 = T1[4'hf:1'h0];
  assign T1 = T44 ? T38 : T2;
  assign T2 = T37 ? T20 : T3;
  assign T3 = T17 ? T11 : twiddle5_4_0_imag;
  assign twiddle5_4_0_imag = T9 + T4;
  assign T4 = {T7, T5};
  assign T5 = $signed(T6) / $signed(22'h100000);
  assign T6 = $signed(1'h0) * $signed(16'hffff);
  assign T7 = T8 ? 31'h7fffffff : 31'h0;
  assign T8 = T5[5'h10:5'h10];
  assign T9 = $signed(T10) / $signed(22'h100000);
  assign T10 = $signed(32'h40000000) * $signed(16'h0);
  assign T11 = {T16, twiddle5_4_1_imag};
  assign twiddle5_4_1_imag = T14 + T12;
  assign T12 = $signed(T13) / $signed(22'h100000);
  assign T13 = $signed(31'h360977fe) * $signed(16'hffff);
  assign T14 = $signed(T15) / $signed(22'h100000);
  assign T15 = $signed(31'h224afc78) * $signed(16'h0);
  assign T16 = twiddle5_4_1_imag[6'h2e:6'h2e];
  assign T17 = T18[1'h0:1'h0];
  assign T18 = T19;
  assign T19 = io_in5[2'h2:1'h0];
  assign T20 = {T36, T21};
  assign T21 = T35 ? twiddle5_4_3_imag : twiddle5_4_2_imag;
  assign twiddle5_4_2_imag = T24 + T22;
  assign T22 = $signed(T23) / $signed(22'h100000);
  assign T23 = $signed(31'h39e8afb9) * $signed(16'hffff);
  assign T24 = {T27, T25};
  assign T25 = $signed(T26) / $signed(22'h100000);
  assign T26 = $signed(30'h24c00837) * $signed(16'h0);
  assign T27 = T25[6'h2d:6'h2d];
  assign twiddle5_4_3_imag = T33 + T28;
  assign T28 = {T31, T29};
  assign T29 = $signed(T30) / $signed(22'h100000);
  assign T30 = $signed(29'h80575ae) * $signed(16'hffff);
  assign T31 = T32 ? 2'h3 : 2'h0;
  assign T32 = T29[6'h2c:6'h2c];
  assign T33 = $signed(T34) / $signed(22'h100000);
  assign T34 = $signed(31'h40813157) * $signed(16'h0);
  assign T35 = T18[1'h0:1'h0];
  assign T36 = T21[6'h2e:6'h2e];
  assign T37 = T18[1'h1:1'h1];
  assign T38 = {T43, twiddle5_4_4_imag};
  assign twiddle5_4_4_imag = T41 + T39;
  assign T39 = $signed(T40) / $signed(22'h100000);
  assign T40 = $signed(31'h4eafe93a) * $signed(16'hffff);
  assign T41 = $signed(T42) / $signed(22'h100000);
  assign T42 = $signed(31'h57347203) * $signed(16'h0);
  assign T43 = twiddle5_4_4_imag[6'h2e:6'h2e];
  assign T44 = T18[2'h2:2'h2];
  assign io_t5_4out_real = T45;
  assign T45 = T46[4'hf:1'h0];
  assign T46 = T87 ? T81 : T47;
  assign T47 = T80 ? T63 : T48;
  assign T48 = T62 ? T56 : twiddle5_4_0_real;
  assign twiddle5_4_0_real = T54 + T49;
  assign T49 = {T52, T50};
  assign T50 = $signed(T51) / $signed(22'h100000);
  assign T51 = $signed(1'h0) * $signed(16'h0);
  assign T52 = T53 ? 31'h7fffffff : 31'h0;
  assign T53 = T50[5'h10:5'h10];
  assign T54 = $signed(T55) / $signed(22'h100000);
  assign T55 = $signed(32'h40000000) * $signed(16'h1);
  assign T56 = {T61, twiddle5_4_1_real};
  assign twiddle5_4_1_real = T59 + T57;
  assign T57 = $signed(T58) / $signed(22'h100000);
  assign T58 = $signed(31'h360977fe) * $signed(16'h0);
  assign T59 = $signed(T60) / $signed(22'h100000);
  assign T60 = $signed(31'h224afc78) * $signed(16'h1);
  assign T61 = twiddle5_4_1_real[6'h2e:6'h2e];
  assign T62 = T18[1'h0:1'h0];
  assign T63 = {T79, T64};
  assign T64 = T78 ? twiddle5_4_3_real : twiddle5_4_2_real;
  assign twiddle5_4_2_real = T67 + T65;
  assign T65 = $signed(T66) / $signed(22'h100000);
  assign T66 = $signed(31'h39e8afb9) * $signed(16'h0);
  assign T67 = {T70, T68};
  assign T68 = $signed(T69) / $signed(22'h100000);
  assign T69 = $signed(30'h24c00837) * $signed(16'h1);
  assign T70 = T68[6'h2d:6'h2d];
  assign twiddle5_4_3_real = T76 + T71;
  assign T71 = {T74, T72};
  assign T72 = $signed(T73) / $signed(22'h100000);
  assign T73 = $signed(29'h80575ae) * $signed(16'h0);
  assign T74 = T75 ? 2'h3 : 2'h0;
  assign T75 = T72[6'h2c:6'h2c];
  assign T76 = $signed(T77) / $signed(22'h100000);
  assign T77 = $signed(31'h40813157) * $signed(16'h1);
  assign T78 = T18[1'h0:1'h0];
  assign T79 = T64[6'h2e:6'h2e];
  assign T80 = T18[1'h1:1'h1];
  assign T81 = {T86, twiddle5_4_4_real};
  assign twiddle5_4_4_real = T84 + T82;
  assign T82 = $signed(T83) / $signed(22'h100000);
  assign T83 = $signed(31'h4eafe93a) * $signed(16'h0);
  assign T84 = $signed(T85) / $signed(22'h100000);
  assign T85 = $signed(31'h57347203) * $signed(16'h1);
  assign T86 = twiddle5_4_4_real[6'h2e:6'h2e];
  assign T87 = T18[2'h2:2'h2];
  assign io_t5_3out_imag = T88;
  assign T88 = T89[4'hf:1'h0];
  assign T89 = T133 ? T124 : T90;
  assign T90 = T123 ? T108 : T91;
  assign T91 = T105 ? T99 : twiddle5_3_0_imag;
  assign twiddle5_3_0_imag = T97 + T92;
  assign T92 = {T95, T93};
  assign T93 = $signed(T94) / $signed(22'h100000);
  assign T94 = $signed(1'h0) * $signed(16'hffff);
  assign T95 = T96 ? 31'h7fffffff : 31'h0;
  assign T96 = T93[5'h10:5'h10];
  assign T97 = $signed(T98) / $signed(22'h100000);
  assign T98 = $signed(32'h40000000) * $signed(16'h0);
  assign T99 = {T104, twiddle5_3_1_imag};
  assign twiddle5_3_1_imag = T102 + T100;
  assign T100 = $signed(T101) / $signed(22'h100000);
  assign T101 = $signed(31'h2bcf9eaa) * $signed(16'hffff);
  assign T102 = $signed(T103) / $signed(22'h100000);
  assign T103 = $signed(31'h2ea76c07) * $signed(16'h0);
  assign T104 = twiddle5_3_1_imag[6'h2e:6'h2e];
  assign T105 = T106[1'h0:1'h0];
  assign T106 = T107;
  assign T107 = io_in5[2'h2:1'h0];
  assign T108 = {T122, T109};
  assign T109 = T121 ? twiddle5_3_3_imag : twiddle5_3_2_imag;
  assign twiddle5_3_2_imag = T112 + T110;
  assign T110 = $signed(T111) / $signed(22'h100000);
  assign T111 = $signed(31'h3fdfab7f) * $signed(16'hffff);
  assign T112 = {T115, T113};
  assign T113 = $signed(T114) / $signed(22'h100000);
  assign T114 = $signed(28'h404c286) * $signed(16'h0);
  assign T115 = T116 ? 3'h7 : 3'h0;
  assign T116 = T113[6'h2b:6'h2b];
  assign twiddle5_3_3_imag = T119 + T117;
  assign T117 = $signed(T118) / $signed(22'h100000);
  assign T118 = $signed(31'h315016c6) * $signed(16'hffff);
  assign T119 = $signed(T120) / $signed(22'h100000);
  assign T120 = $signed(31'h57347203) * $signed(16'h0);
  assign T121 = T106[1'h0:1'h0];
  assign T122 = T109[6'h2e:6'h2e];
  assign T123 = T106[1'h1:1'h1];
  assign T124 = {T132, twiddle5_3_4_imag};
  assign twiddle5_3_4_imag = T130 + T125;
  assign T125 = {T128, T126};
  assign T126 = $signed(T127) / $signed(22'h100000);
  assign T127 = $signed(29'h80575ae) * $signed(16'hffff);
  assign T128 = T129 ? 2'h3 : 2'h0;
  assign T129 = T126[6'h2c:6'h2c];
  assign T130 = $signed(T131) / $signed(22'h100000);
  assign T131 = $signed(31'h40813157) * $signed(16'h0);
  assign T132 = twiddle5_3_4_imag[6'h2e:6'h2e];
  assign T133 = T106[2'h2:2'h2];
  assign io_t5_3out_real = T134;
  assign T134 = T135[4'hf:1'h0];
  assign T135 = T177 ? T168 : T136;
  assign T136 = T167 ? T152 : T137;
  assign T137 = T151 ? T145 : twiddle5_3_0_real;
  assign twiddle5_3_0_real = T143 + T138;
  assign T138 = {T141, T139};
  assign T139 = $signed(T140) / $signed(22'h100000);
  assign T140 = $signed(1'h0) * $signed(16'h0);
  assign T141 = T142 ? 31'h7fffffff : 31'h0;
  assign T142 = T139[5'h10:5'h10];
  assign T143 = $signed(T144) / $signed(22'h100000);
  assign T144 = $signed(32'h40000000) * $signed(16'h1);
  assign T145 = {T150, twiddle5_3_1_real};
  assign twiddle5_3_1_real = T148 + T146;
  assign T146 = $signed(T147) / $signed(22'h100000);
  assign T147 = $signed(31'h2bcf9eaa) * $signed(16'h0);
  assign T148 = $signed(T149) / $signed(22'h100000);
  assign T149 = $signed(31'h2ea76c07) * $signed(16'h1);
  assign T150 = twiddle5_3_1_real[6'h2e:6'h2e];
  assign T151 = T106[1'h0:1'h0];
  assign T152 = {T166, T153};
  assign T153 = T165 ? twiddle5_3_3_real : twiddle5_3_2_real;
  assign twiddle5_3_2_real = T156 + T154;
  assign T154 = $signed(T155) / $signed(22'h100000);
  assign T155 = $signed(31'h3fdfab7f) * $signed(16'h0);
  assign T156 = {T159, T157};
  assign T157 = $signed(T158) / $signed(22'h100000);
  assign T158 = $signed(28'h404c286) * $signed(16'h1);
  assign T159 = T160 ? 3'h7 : 3'h0;
  assign T160 = T157[6'h2b:6'h2b];
  assign twiddle5_3_3_real = T163 + T161;
  assign T161 = $signed(T162) / $signed(22'h100000);
  assign T162 = $signed(31'h315016c6) * $signed(16'h0);
  assign T163 = $signed(T164) / $signed(22'h100000);
  assign T164 = $signed(31'h57347203) * $signed(16'h1);
  assign T165 = T106[1'h0:1'h0];
  assign T166 = T153[6'h2e:6'h2e];
  assign T167 = T106[1'h1:1'h1];
  assign T168 = {T176, twiddle5_3_4_real};
  assign twiddle5_3_4_real = T174 + T169;
  assign T169 = {T172, T170};
  assign T170 = $signed(T171) / $signed(22'h100000);
  assign T171 = $signed(29'h80575ae) * $signed(16'h0);
  assign T172 = T173 ? 2'h3 : 2'h0;
  assign T173 = T170[6'h2c:6'h2c];
  assign T174 = $signed(T175) / $signed(22'h100000);
  assign T175 = $signed(31'h40813157) * $signed(16'h1);
  assign T176 = twiddle5_3_4_real[6'h2e:6'h2e];
  assign T177 = T106[2'h2:2'h2];
  assign io_t5_2out_imag = T178;
  assign T178 = T179[4'hf:1'h0];
  assign T179 = T224 ? T216 : T180;
  assign T180 = T215 ? T200 : T181;
  assign T181 = T197 ? T189 : twiddle5_2_0_imag;
  assign twiddle5_2_0_imag = T187 + T182;
  assign T182 = {T185, T183};
  assign T183 = $signed(T184) / $signed(22'h100000);
  assign T184 = $signed(1'h0) * $signed(16'hffff);
  assign T185 = T186 ? 31'h7fffffff : 31'h0;
  assign T186 = T183[5'h10:5'h10];
  assign T187 = $signed(T188) / $signed(22'h100000);
  assign T188 = $signed(32'h40000000) * $signed(16'h0);
  assign T189 = {T196, twiddle5_2_1_imag};
  assign twiddle5_2_1_imag = T194 + T190;
  assign T190 = {T193, T191};
  assign T191 = $signed(T192) / $signed(22'h100000);
  assign T192 = $signed(30'h1ed50d5c) * $signed(16'hffff);
  assign T193 = T191[6'h2d:6'h2d];
  assign T194 = $signed(T195) / $signed(22'h100000);
  assign T195 = $signed(31'h3815689d) * $signed(16'h0);
  assign T196 = twiddle5_2_1_imag[6'h2e:6'h2e];
  assign T197 = T198[1'h0:1'h0];
  assign T198 = T199;
  assign T199 = io_in5[2'h2:1'h0];
  assign T200 = {T214, T201};
  assign T201 = T213 ? twiddle5_2_3_imag : twiddle5_2_2_imag;
  assign twiddle5_2_2_imag = T204 + T202;
  assign T202 = $signed(T203) / $signed(22'h100000);
  assign T203 = $signed(31'h360977fe) * $signed(16'hffff);
  assign T204 = $signed(T205) / $signed(22'h100000);
  assign T205 = $signed(31'h224afc78) * $signed(16'h0);
  assign twiddle5_2_3_imag = T208 + T206;
  assign T206 = $signed(T207) / $signed(22'h100000);
  assign T207 = $signed(31'h3fdfab7f) * $signed(16'hffff);
  assign T208 = {T211, T209};
  assign T209 = $signed(T210) / $signed(22'h100000);
  assign T210 = $signed(28'h404c286) * $signed(16'h0);
  assign T211 = T212 ? 3'h7 : 3'h0;
  assign T212 = T209[6'h2b:6'h2b];
  assign T213 = T198[1'h0:1'h0];
  assign T214 = T201[6'h2e:6'h2e];
  assign T215 = T198[1'h1:1'h1];
  assign T216 = {T223, twiddle5_2_4_imag};
  assign twiddle5_2_4_imag = T219 + T217;
  assign T217 = $signed(T218) / $signed(22'h100000);
  assign T218 = $signed(31'h39e8afb9) * $signed(16'hffff);
  assign T219 = {T222, T220};
  assign T220 = $signed(T221) / $signed(22'h100000);
  assign T221 = $signed(30'h24c00837) * $signed(16'h0);
  assign T222 = T220[6'h2d:6'h2d];
  assign T223 = twiddle5_2_4_imag[6'h2e:6'h2e];
  assign T224 = T198[2'h2:2'h2];
  assign io_t5_2out_real = T225;
  assign T225 = T226[4'hf:1'h0];
  assign T226 = T269 ? T261 : T227;
  assign T227 = T260 ? T245 : T228;
  assign T228 = T244 ? T236 : twiddle5_2_0_real;
  assign twiddle5_2_0_real = T234 + T229;
  assign T229 = {T232, T230};
  assign T230 = $signed(T231) / $signed(22'h100000);
  assign T231 = $signed(1'h0) * $signed(16'h0);
  assign T232 = T233 ? 31'h7fffffff : 31'h0;
  assign T233 = T230[5'h10:5'h10];
  assign T234 = $signed(T235) / $signed(22'h100000);
  assign T235 = $signed(32'h40000000) * $signed(16'h1);
  assign T236 = {T243, twiddle5_2_1_real};
  assign twiddle5_2_1_real = T241 + T237;
  assign T237 = {T240, T238};
  assign T238 = $signed(T239) / $signed(22'h100000);
  assign T239 = $signed(30'h1ed50d5c) * $signed(16'h0);
  assign T240 = T238[6'h2d:6'h2d];
  assign T241 = $signed(T242) / $signed(22'h100000);
  assign T242 = $signed(31'h3815689d) * $signed(16'h1);
  assign T243 = twiddle5_2_1_real[6'h2e:6'h2e];
  assign T244 = T198[1'h0:1'h0];
  assign T245 = {T259, T246};
  assign T246 = T258 ? twiddle5_2_3_real : twiddle5_2_2_real;
  assign twiddle5_2_2_real = T249 + T247;
  assign T247 = $signed(T248) / $signed(22'h100000);
  assign T248 = $signed(31'h360977fe) * $signed(16'h0);
  assign T249 = $signed(T250) / $signed(22'h100000);
  assign T250 = $signed(31'h224afc78) * $signed(16'h1);
  assign twiddle5_2_3_real = T253 + T251;
  assign T251 = $signed(T252) / $signed(22'h100000);
  assign T252 = $signed(31'h3fdfab7f) * $signed(16'h0);
  assign T253 = {T256, T254};
  assign T254 = $signed(T255) / $signed(22'h100000);
  assign T255 = $signed(28'h404c286) * $signed(16'h1);
  assign T256 = T257 ? 3'h7 : 3'h0;
  assign T257 = T254[6'h2b:6'h2b];
  assign T258 = T198[1'h0:1'h0];
  assign T259 = T246[6'h2e:6'h2e];
  assign T260 = T198[1'h1:1'h1];
  assign T261 = {T268, twiddle5_2_4_real};
  assign twiddle5_2_4_real = T264 + T262;
  assign T262 = $signed(T263) / $signed(22'h100000);
  assign T263 = $signed(31'h39e8afb9) * $signed(16'h0);
  assign T264 = {T267, T265};
  assign T265 = $signed(T266) / $signed(22'h100000);
  assign T266 = $signed(30'h24c00837) * $signed(16'h1);
  assign T267 = T265[6'h2d:6'h2d];
  assign T268 = twiddle5_2_4_real[6'h2e:6'h2e];
  assign T269 = T198[2'h2:2'h2];
  assign io_t5_1out_imag = T270;
  assign T270 = T271[4'hf:1'h0];
  assign T271 = T314 ? T308 : T272;
  assign T272 = T307 ? T293 : T273;
  assign T273 = T290 ? T281 : twiddle5_1_0_imag;
  assign twiddle5_1_0_imag = T279 + T274;
  assign T274 = {T277, T275};
  assign T275 = $signed(T276) / $signed(22'h100000);
  assign T276 = $signed(1'h0) * $signed(16'hffff);
  assign T277 = T278 ? 31'h7fffffff : 31'h0;
  assign T278 = T275[5'h10:5'h10];
  assign T279 = $signed(T280) / $signed(22'h100000);
  assign T280 = $signed(32'h40000000) * $signed(16'h0);
  assign T281 = {T289, twiddle5_1_1_imag};
  assign twiddle5_1_1_imag = T287 + T282;
  assign T282 = {T285, T283};
  assign T283 = $signed(T284) / $signed(22'h100000);
  assign T284 = $signed(29'hfea88fd) * $signed(16'hffff);
  assign T285 = T286 ? 2'h3 : 2'h0;
  assign T286 = T283[6'h2c:6'h2c];
  assign T287 = $signed(T288) / $signed(22'h100000);
  assign T288 = $signed(31'h3dfd443a) * $signed(16'h0);
  assign T289 = twiddle5_1_1_imag[6'h2e:6'h2e];
  assign T290 = T291[1'h0:1'h0];
  assign T291 = T292;
  assign T292 = io_in5[2'h2:1'h0];
  assign T293 = {T306, T294};
  assign T294 = T305 ? twiddle5_1_3_imag : twiddle5_1_2_imag;
  assign twiddle5_1_2_imag = T299 + T295;
  assign T295 = {T298, T296};
  assign T296 = $signed(T297) / $signed(22'h100000);
  assign T297 = $signed(30'h1ed50d5c) * $signed(16'hffff);
  assign T298 = T296[6'h2d:6'h2d];
  assign T299 = $signed(T300) / $signed(22'h100000);
  assign T300 = $signed(31'h3815689d) * $signed(16'h0);
  assign twiddle5_1_3_imag = T303 + T301;
  assign T301 = $signed(T302) / $signed(22'h100000);
  assign T302 = $signed(31'h2bcf9eaa) * $signed(16'hffff);
  assign T303 = $signed(T304) / $signed(22'h100000);
  assign T304 = $signed(31'h2ea76c07) * $signed(16'h0);
  assign T305 = T291[1'h0:1'h0];
  assign T306 = T294[6'h2e:6'h2e];
  assign T307 = T291[1'h1:1'h1];
  assign T308 = {T313, twiddle5_1_4_imag};
  assign twiddle5_1_4_imag = T311 + T309;
  assign T309 = $signed(T310) / $signed(22'h100000);
  assign T310 = $signed(31'h360977fe) * $signed(16'hffff);
  assign T311 = $signed(T312) / $signed(22'h100000);
  assign T312 = $signed(31'h224afc78) * $signed(16'h0);
  assign T313 = twiddle5_1_4_imag[6'h2e:6'h2e];
  assign T314 = T291[2'h2:2'h2];
  assign io_t5_1out_real = T315;
  assign T315 = T316[4'hf:1'h0];
  assign T316 = T357 ? T351 : T317;
  assign T317 = T350 ? T336 : T318;
  assign T318 = T335 ? T326 : twiddle5_1_0_real;
  assign twiddle5_1_0_real = T324 + T319;
  assign T319 = {T322, T320};
  assign T320 = $signed(T321) / $signed(22'h100000);
  assign T321 = $signed(1'h0) * $signed(16'h0);
  assign T322 = T323 ? 31'h7fffffff : 31'h0;
  assign T323 = T320[5'h10:5'h10];
  assign T324 = $signed(T325) / $signed(22'h100000);
  assign T325 = $signed(32'h40000000) * $signed(16'h1);
  assign T326 = {T334, twiddle5_1_1_real};
  assign twiddle5_1_1_real = T332 + T327;
  assign T327 = {T330, T328};
  assign T328 = $signed(T329) / $signed(22'h100000);
  assign T329 = $signed(29'hfea88fd) * $signed(16'h0);
  assign T330 = T331 ? 2'h3 : 2'h0;
  assign T331 = T328[6'h2c:6'h2c];
  assign T332 = $signed(T333) / $signed(22'h100000);
  assign T333 = $signed(31'h3dfd443a) * $signed(16'h1);
  assign T334 = twiddle5_1_1_real[6'h2e:6'h2e];
  assign T335 = T291[1'h0:1'h0];
  assign T336 = {T349, T337};
  assign T337 = T348 ? twiddle5_1_3_real : twiddle5_1_2_real;
  assign twiddle5_1_2_real = T342 + T338;
  assign T338 = {T341, T339};
  assign T339 = $signed(T340) / $signed(22'h100000);
  assign T340 = $signed(30'h1ed50d5c) * $signed(16'h0);
  assign T341 = T339[6'h2d:6'h2d];
  assign T342 = $signed(T343) / $signed(22'h100000);
  assign T343 = $signed(31'h3815689d) * $signed(16'h1);
  assign twiddle5_1_3_real = T346 + T344;
  assign T344 = $signed(T345) / $signed(22'h100000);
  assign T345 = $signed(31'h2bcf9eaa) * $signed(16'h0);
  assign T346 = $signed(T347) / $signed(22'h100000);
  assign T347 = $signed(31'h2ea76c07) * $signed(16'h1);
  assign T348 = T291[1'h0:1'h0];
  assign T349 = T337[6'h2e:6'h2e];
  assign T350 = T291[1'h1:1'h1];
  assign T351 = {T356, twiddle5_1_4_real};
  assign twiddle5_1_4_real = T354 + T352;
  assign T352 = $signed(T353) / $signed(22'h100000);
  assign T353 = $signed(31'h360977fe) * $signed(16'h0);
  assign T354 = $signed(T355) / $signed(22'h100000);
  assign T355 = $signed(31'h224afc78) * $signed(16'h1);
  assign T356 = twiddle5_1_4_real[6'h2e:6'h2e];
  assign T357 = T291[2'h2:2'h2];
  assign io_t3_2out_imag = T358;
  assign T358 = T359[4'hf:1'h0];
  assign T359 = T985 ? T867 : T360;
  assign T360 = T866 ? T618 : T361;
  assign T361 = T617 ? T493 : T362;
  assign T362 = T492 ? T438 : T363;
  assign T363 = T437 ? T404 : T364;
  assign T364 = T403 ? T385 : T365;
  assign T365 = T382 ? T373 : twiddle3_2_0_imag;
  assign twiddle3_2_0_imag = T371 + T366;
  assign T366 = {T369, T367};
  assign T367 = $signed(T368) / $signed(22'h100000);
  assign T368 = $signed(1'h0) * $signed(16'hffff);
  assign T369 = T370 ? 31'h7fffffff : 31'h0;
  assign T370 = T367[5'h10:5'h10];
  assign T371 = $signed(T372) / $signed(22'h100000);
  assign T372 = $signed(32'h40000000) * $signed(16'h0);
  assign T373 = {T381, twiddle3_2_1_imag};
  assign twiddle3_2_1_imag = T379 + T374;
  assign T374 = {T377, T375};
  assign T375 = $signed(T376) / $signed(22'h100000);
  assign T376 = $signed(27'h34ee54e) * $signed(16'hffff);
  assign T377 = T378 ? 4'hf : 4'h0;
  assign T378 = T375[6'h2a:6'h2a];
  assign T379 = $signed(T380) / $signed(22'h100000);
  assign T380 = $signed(31'h3fea18df) * $signed(16'h0);
  assign T381 = twiddle3_2_1_imag[6'h2e:6'h2e];
  assign T382 = T383[1'h0:1'h0];
  assign T383 = T384;
  assign T384 = io_in3[3'h6:1'h0];
  assign T385 = {T402, T386};
  assign T386 = T401 ? twiddle3_2_3_imag : twiddle3_2_2_imag;
  assign twiddle3_2_2_imag = T392 + T387;
  assign T387 = {T390, T388};
  assign T388 = $signed(T389) / $signed(22'h100000);
  assign T389 = $signed(28'h69b86f1) * $signed(16'hffff);
  assign T390 = T391 ? 3'h7 : 3'h0;
  assign T391 = T388[6'h2b:6'h2b];
  assign T392 = $signed(T393) / $signed(22'h100000);
  assign T393 = $signed(31'h3fa8727d) * $signed(16'h0);
  assign twiddle3_2_3_imag = T399 + T394;
  assign T394 = {T397, T395};
  assign T395 = $signed(T396) / $signed(22'h100000);
  assign T396 = $signed(29'h9e3a2ca) * $signed(16'hffff);
  assign T397 = T398 ? 2'h3 : 2'h0;
  assign T398 = T395[6'h2c:6'h2c];
  assign T399 = $signed(T400) / $signed(22'h100000);
  assign T400 = $signed(31'h3f3b39c7) * $signed(16'h0);
  assign T401 = T383[1'h0:1'h0];
  assign T402 = T386[6'h2e:6'h2e];
  assign T403 = T383[1'h1:1'h1];
  assign T404 = {T436, T405};
  assign T405 = T435 ? T421 : T406;
  assign T406 = T420 ? twiddle3_2_5_imag : twiddle3_2_4_imag;
  assign twiddle3_2_4_imag = T412 + T407;
  assign T407 = {T410, T408};
  assign T408 = $signed(T409) / $signed(22'h100000);
  assign T409 = $signed(29'hd24f9d3) * $signed(16'hffff);
  assign T410 = T411 ? 2'h3 : 2'h0;
  assign T411 = T408[6'h2c:6'h2c];
  assign T412 = $signed(T413) / $signed(22'h100000);
  assign T413 = $signed(31'h3ea2b980) * $signed(16'h0);
  assign twiddle3_2_5_imag = T418 + T414;
  assign T414 = {T417, T415};
  assign T415 = $signed(T416) / $signed(22'h100000);
  assign T416 = $signed(30'h105d51a8) * $signed(16'hffff);
  assign T417 = T415[6'h2d:6'h2d];
  assign T418 = $signed(T419) / $signed(22'h100000);
  assign T419 = $signed(31'h3ddf5a09) * $signed(16'h0);
  assign T420 = T383[1'h0:1'h0];
  assign T421 = T434 ? twiddle3_2_7_imag : twiddle3_2_6_imag;
  assign twiddle3_2_6_imag = T426 + T422;
  assign T422 = {T425, T423};
  assign T423 = $signed(T424) / $signed(22'h100000);
  assign T424 = $signed(30'h138a760d) * $signed(16'hffff);
  assign T425 = T423[6'h2d:6'h2d];
  assign T426 = $signed(T427) / $signed(22'h100000);
  assign T427 = $signed(31'h3cf1a11d) * $signed(16'h0);
  assign twiddle3_2_7_imag = T432 + T428;
  assign T428 = {T431, T429};
  assign T429 = $signed(T430) / $signed(22'h100000);
  assign T430 = $signed(30'h16aa3a72) * $signed(16'hffff);
  assign T431 = T429[6'h2d:6'h2d];
  assign T432 = $signed(T433) / $signed(22'h100000);
  assign T433 = $signed(31'h3bda3171) * $signed(16'h0);
  assign T434 = T383[1'h0:1'h0];
  assign T435 = T383[1'h1:1'h1];
  assign T436 = T405[6'h2e:6'h2e];
  assign T437 = T383[2'h2:2'h2];
  assign T438 = {T491, T439};
  assign T439 = T490 ? T468 : T440;
  assign T440 = T467 ? T455 : T441;
  assign T441 = T454 ? twiddle3_2_9_imag : twiddle3_2_8_imag;
  assign twiddle3_2_8_imag = T446 + T442;
  assign T442 = {T445, T443};
  assign T443 = $signed(T444) / $signed(22'h100000);
  assign T444 = $signed(30'h19ba7b6c) * $signed(16'hffff);
  assign T445 = T443[6'h2d:6'h2d];
  assign T446 = $signed(T447) / $signed(22'h100000);
  assign T447 = $signed(31'h3a99ca4a) * $signed(16'h0);
  assign twiddle3_2_9_imag = T452 + T448;
  assign T448 = {T451, T449};
  assign T449 = $signed(T450) / $signed(22'h100000);
  assign T450 = $signed(30'h1cb92032) * $signed(16'hffff);
  assign T451 = T449[6'h2d:6'h2d];
  assign T452 = $signed(T453) / $signed(22'h100000);
  assign T453 = $signed(31'h393146f5) * $signed(16'h0);
  assign T454 = T383[1'h0:1'h0];
  assign T455 = T466 ? twiddle3_2_11_imag : twiddle3_2_10_imag;
  assign twiddle3_2_10_imag = T460 + T456;
  assign T456 = {T459, T457};
  assign T457 = $signed(T458) / $signed(22'h100000);
  assign T458 = $signed(30'h1fa41c05) * $signed(16'hffff);
  assign T459 = T457[6'h2d:6'h2d];
  assign T460 = $signed(T461) / $signed(22'h100000);
  assign T461 = $signed(31'h37a19e34) * $signed(16'h0);
  assign twiddle3_2_11_imag = T464 + T462;
  assign T462 = $signed(T463) / $signed(22'h100000);
  assign T463 = $signed(31'h22796f9d) * $signed(16'hffff);
  assign T464 = $signed(T465) / $signed(22'h100000);
  assign T465 = $signed(31'h35ebe194) * $signed(16'h0);
  assign T466 = T383[1'h0:1'h0];
  assign T467 = T383[1'h1:1'h1];
  assign T468 = T489 ? T479 : T469;
  assign T469 = T478 ? twiddle3_2_13_imag : twiddle3_2_12_imag;
  assign twiddle3_2_12_imag = T472 + T470;
  assign T470 = $signed(T471) / $signed(22'h100000);
  assign T471 = $signed(31'h25372a85) * $signed(16'hffff);
  assign T472 = $signed(T473) / $signed(22'h100000);
  assign T473 = $signed(31'h34113cb3) * $signed(16'h0);
  assign twiddle3_2_13_imag = T476 + T474;
  assign T474 = $signed(T475) / $signed(22'h100000);
  assign T475 = $signed(31'h27db6c6d) * $signed(16'hffff);
  assign T476 = $signed(T477) / $signed(22'h100000);
  assign T477 = $signed(31'h3212f472) * $signed(16'h0);
  assign T478 = T383[1'h0:1'h0];
  assign T479 = T488 ? twiddle3_2_15_imag : twiddle3_2_14_imag;
  assign twiddle3_2_14_imag = T482 + T480;
  assign T480 = $signed(T481) / $signed(22'h100000);
  assign T481 = $signed(31'h2a646676) * $signed(16'hffff);
  assign T482 = $signed(T483) / $signed(22'h100000);
  assign T483 = $signed(31'h2ff26615) * $signed(16'h0);
  assign twiddle3_2_15_imag = T486 + T484;
  assign T484 = $signed(T485) / $signed(22'h100000);
  assign T485 = $signed(31'h2cd05c6c) * $signed(16'hffff);
  assign T486 = $signed(T487) / $signed(22'h100000);
  assign T487 = $signed(31'h2db10657) * $signed(16'h0);
  assign T488 = T383[1'h0:1'h0];
  assign T489 = T383[1'h1:1'h1];
  assign T490 = T383[2'h2:2'h2];
  assign T491 = T439[6'h2e:6'h2e];
  assign T492 = T383[2'h3:2'h3];
  assign T493 = {T616, T494};
  assign T494 = T615 ? T547 : T495;
  assign T495 = T546 ? T518 : T496;
  assign T496 = T517 ? T507 : T497;
  assign T497 = T506 ? twiddle3_2_17_imag : twiddle3_2_16_imag;
  assign twiddle3_2_16_imag = T500 + T498;
  assign T498 = $signed(T499) / $signed(22'h100000);
  assign T499 = $signed(31'h2f1da5f8) * $signed(16'hffff);
  assign T500 = $signed(T501) / $signed(22'h100000);
  assign T501 = $signed(31'h2b506069) * $signed(16'h0);
  assign twiddle3_2_17_imag = T504 + T502;
  assign T502 = $signed(T503) / $signed(22'h100000);
  assign T503 = $signed(31'h314aafc2) * $signed(16'hffff);
  assign T504 = $signed(T505) / $signed(22'h100000);
  assign T505 = $signed(31'h28d214e4) * $signed(16'h0);
  assign T506 = T383[1'h0:1'h0];
  assign T507 = T516 ? twiddle3_2_19_imag : twiddle3_2_18_imag;
  assign twiddle3_2_18_imag = T510 + T508;
  assign T508 = $signed(T509) / $signed(22'h100000);
  assign T509 = $signed(31'h3355fc84) * $signed(16'hffff);
  assign T510 = $signed(T511) / $signed(22'h100000);
  assign T511 = $signed(31'h2637d8ab) * $signed(16'h0);
  assign twiddle3_2_19_imag = T514 + T512;
  assign T512 = $signed(T513) / $signed(22'h100000);
  assign T513 = $signed(31'h353e260f) * $signed(16'hffff);
  assign T514 = $signed(T515) / $signed(22'h100000);
  assign T515 = $signed(31'h238373c3) * $signed(16'h0);
  assign T516 = T383[1'h0:1'h0];
  assign T517 = T383[1'h1:1'h1];
  assign T518 = T545 ? T531 : T519;
  assign T519 = T530 ? twiddle3_2_21_imag : twiddle3_2_20_imag;
  assign twiddle3_2_20_imag = T522 + T520;
  assign T520 = $signed(T521) / $signed(22'h100000);
  assign T521 = $signed(31'h3701de44) * $signed(16'hffff);
  assign T522 = $signed(T523) / $signed(22'h100000);
  assign T523 = $signed(31'h20b6c016) * $signed(16'h0);
  assign twiddle3_2_21_imag = T526 + T524;
  assign T524 = $signed(T525) / $signed(22'h100000);
  assign T525 = $signed(31'h389feff1) * $signed(16'hffff);
  assign T526 = {T529, T527};
  assign T527 = $signed(T528) / $signed(22'h100000);
  assign T528 = $signed(30'h1dd3a832) * $signed(16'h0);
  assign T529 = T527[6'h2d:6'h2d];
  assign T530 = T383[1'h0:1'h0];
  assign T531 = T544 ? twiddle3_2_23_imag : twiddle3_2_22_imag;
  assign twiddle3_2_22_imag = T534 + T532;
  assign T532 = $signed(T533) / $signed(22'h100000);
  assign T533 = $signed(31'h3a173fae) * $signed(16'hffff);
  assign T534 = {T537, T535};
  assign T535 = $signed(T536) / $signed(22'h100000);
  assign T536 = $signed(30'h1adc25fb) * $signed(16'h0);
  assign T537 = T535[6'h2d:6'h2d];
  assign twiddle3_2_23_imag = T540 + T538;
  assign T538 = $signed(T539) / $signed(22'h100000);
  assign T539 = $signed(31'h3b66cc97) * $signed(16'hffff);
  assign T540 = {T543, T541};
  assign T541 = $signed(T542) / $signed(22'h100000);
  assign T542 = $signed(30'h17d2414a) * $signed(16'h0);
  assign T543 = T541[6'h2d:6'h2d];
  assign T544 = T383[1'h0:1'h0];
  assign T545 = T383[1'h1:1'h1];
  assign T546 = T383[2'h2:2'h2];
  assign T547 = T614 ? T580 : T548;
  assign T548 = T579 ? T563 : T549;
  assign T549 = T562 ? twiddle3_2_25_imag : twiddle3_2_24_imag;
  assign twiddle3_2_24_imag = T552 + T550;
  assign T550 = $signed(T551) / $signed(22'h100000);
  assign T551 = $signed(31'h3c8db0ff) * $signed(16'hffff);
  assign T552 = {T555, T553};
  assign T553 = $signed(T554) / $signed(22'h100000);
  assign T554 = $signed(30'h14b80e91) * $signed(16'h0);
  assign T555 = T553[6'h2d:6'h2d];
  assign twiddle3_2_25_imag = T558 + T556;
  assign T556 = $signed(T557) / $signed(22'h100000);
  assign T557 = $signed(31'h3d8b2310) * $signed(16'hffff);
  assign T558 = {T561, T559};
  assign T559 = $signed(T560) / $signed(22'h100000);
  assign T560 = $signed(30'h118fad69) * $signed(16'h0);
  assign T561 = T559[6'h2d:6'h2d];
  assign T562 = T383[1'h0:1'h0];
  assign T563 = T578 ? twiddle3_2_27_imag : twiddle3_2_26_imag;
  assign twiddle3_2_26_imag = T566 + T564;
  assign T564 = $signed(T565) / $signed(22'h100000);
  assign T565 = $signed(31'h3e5e754f) * $signed(16'hffff);
  assign T566 = {T569, T567};
  assign T567 = $signed(T568) / $signed(22'h100000);
  assign T568 = $signed(29'he5b4720) * $signed(16'h0);
  assign T569 = T570 ? 2'h3 : 2'h0;
  assign T570 = T567[6'h2c:6'h2c];
  assign twiddle3_2_27_imag = T573 + T571;
  assign T571 = $signed(T572) / $signed(22'h100000);
  assign T572 = $signed(31'h3f071719) * $signed(16'hffff);
  assign T573 = {T576, T574};
  assign T574 = $signed(T575) / $signed(22'h100000);
  assign T575 = $signed(29'hb1d0d3f) * $signed(16'h0);
  assign T576 = T577 ? 2'h3 : 2'h0;
  assign T577 = T574[6'h2c:6'h2c];
  assign T578 = T383[1'h0:1'h0];
  assign T579 = T383[1'h1:1'h1];
  assign T580 = T613 ? T597 : T581;
  assign T581 = T596 ? twiddle3_2_29_imag : twiddle3_2_28_imag;
  assign twiddle3_2_28_imag = T584 + T582;
  assign T582 = $signed(T583) / $signed(22'h100000);
  assign T583 = $signed(31'h3f849500) * $signed(16'hffff);
  assign T584 = {T587, T585};
  assign T585 = $signed(T586) / $signed(22'h100000);
  assign T586 = $signed(28'h7d73808) * $signed(16'h0);
  assign T587 = T588 ? 3'h7 : 3'h0;
  assign T588 = T585[6'h2b:6'h2b];
  assign twiddle3_2_29_imag = T591 + T589;
  assign T589 = $signed(T590) / $signed(22'h100000);
  assign T590 = $signed(31'h3fd69921) * $signed(16'hffff);
  assign T591 = {T594, T592};
  assign T592 = $signed(T593) / $signed(22'h100000);
  assign T593 = $signed(28'h48c04f3) * $signed(16'h0);
  assign T594 = T595 ? 3'h7 : 3'h0;
  assign T595 = T592[6'h2b:6'h2b];
  assign T596 = T383[1'h0:1'h0];
  assign T597 = T612 ? twiddle3_2_31_imag : twiddle3_2_30_imag;
  assign twiddle3_2_30_imag = T600 + T598;
  assign T598 = $signed(T599) / $signed(22'h100000);
  assign T599 = $signed(31'h3ffceb58) * $signed(16'hffff);
  assign T600 = {T603, T601};
  assign T601 = $signed(T602) / $signed(22'h100000);
  assign T602 = $signed(26'h13db523) * $signed(16'h0);
  assign T603 = T604 ? 5'h1f : 5'h0;
  assign T604 = T601[6'h29:6'h29];
  assign twiddle3_2_31_imag = T607 + T605;
  assign T605 = $signed(T606) / $signed(22'h100000);
  assign T606 = $signed(31'h3ff7716b) * $signed(16'hffff);
  assign T607 = {T610, T608};
  assign T608 = $signed(T609) / $signed(22'h100000);
  assign T609 = $signed(27'h5ee8bdf) * $signed(16'h0);
  assign T610 = T611 ? 4'hf : 4'h0;
  assign T611 = T608[6'h2a:6'h2a];
  assign T612 = T383[1'h0:1'h0];
  assign T613 = T383[1'h1:1'h1];
  assign T614 = T383[2'h2:2'h2];
  assign T615 = T383[2'h3:2'h3];
  assign T616 = T494[6'h2e:6'h2e];
  assign T617 = T383[3'h4:3'h4];
  assign T618 = {T865, T619};
  assign T619 = T864 ? T736 : T620;
  assign T620 = T735 ? T687 : T621;
  assign T621 = T686 ? T656 : T622;
  assign T622 = T655 ? T639 : T623;
  assign T623 = T638 ? twiddle3_2_33_imag : twiddle3_2_32_imag;
  assign twiddle3_2_32_imag = T626 + T624;
  assign T624 = $signed(T625) / $signed(22'h100000);
  assign T625 = $signed(31'h3fc62f18) * $signed(16'hffff);
  assign T626 = {T629, T627};
  assign T627 = $signed(T628) / $signed(22'h100000);
  assign T628 = $signed(28'haa0ccff) * $signed(16'h0);
  assign T629 = T630 ? 3'h7 : 3'h0;
  assign T630 = T627[6'h2b:6'h2b];
  assign twiddle3_2_33_imag = T633 + T631;
  assign T631 = $signed(T632) / $signed(22'h100000);
  assign T632 = $signed(31'h3f694618) * $signed(16'hffff);
  assign T633 = {T636, T634};
  assign T634 = $signed(T635) / $signed(22'h100000);
  assign T635 = $signed(29'h1756bb64) * $signed(16'h0);
  assign T636 = T637 ? 2'h3 : 2'h0;
  assign T637 = T634[6'h2c:6'h2c];
  assign T638 = T383[1'h0:1'h0];
  assign T639 = T654 ? twiddle3_2_35_imag : twiddle3_2_34_imag;
  assign twiddle3_2_34_imag = T642 + T640;
  assign T640 = $signed(T641) / $signed(22'h100000);
  assign T641 = $signed(31'h3ee0f602) * $signed(16'hffff);
  assign T642 = {T645, T643};
  assign T643 = $signed(T644) / $signed(22'h100000);
  assign T644 = $signed(29'h1412976d) * $signed(16'h0);
  assign T645 = T646 ? 2'h3 : 2'h0;
  assign T646 = T643[6'h2c:6'h2c];
  assign twiddle3_2_35_imag = T649 + T647;
  assign T647 = $signed(T648) / $signed(22'h100000);
  assign T648 = $signed(31'h3e2d9c23) * $signed(16'hffff);
  assign T649 = {T652, T650};
  assign T650 = $signed(T651) / $signed(22'h100000);
  assign T651 = $signed(29'h10d69d68) * $signed(16'h0);
  assign T652 = T653 ? 2'h3 : 2'h0;
  assign T653 = T650[6'h2c:6'h2c];
  assign T654 = T383[1'h0:1'h0];
  assign T655 = T383[1'h1:1'h1];
  assign T656 = T685 ? T671 : T657;
  assign T657 = T670 ? twiddle3_2_37_imag : twiddle3_2_36_imag;
  assign twiddle3_2_36_imag = T660 + T658;
  assign T658 = $signed(T659) / $signed(22'h100000);
  assign T659 = $signed(31'h3d4fb33e) * $signed(16'hffff);
  assign T660 = {T663, T661};
  assign T661 = $signed(T662) / $signed(22'h100000);
  assign T662 = $signed(30'h2da5040e) * $signed(16'h0);
  assign T663 = T661[6'h2d:6'h2d];
  assign twiddle3_2_37_imag = T666 + T664;
  assign T664 = $signed(T665) / $signed(22'h100000);
  assign T665 = $signed(31'h3c47d336) * $signed(16'hffff);
  assign T666 = {T669, T667};
  assign T667 = $signed(T668) / $signed(22'h100000);
  assign T668 = $signed(30'h2a7ffafd) * $signed(16'h0);
  assign T669 = T667[6'h2d:6'h2d];
  assign T670 = T383[1'h0:1'h0];
  assign T671 = T684 ? twiddle3_2_39_imag : twiddle3_2_38_imag;
  assign twiddle3_2_38_imag = T674 + T672;
  assign T672 = $signed(T673) / $signed(22'h100000);
  assign T673 = $signed(31'h3b16b0a8) * $signed(16'hffff);
  assign T674 = {T677, T675};
  assign T675 = $signed(T676) / $signed(22'h100000);
  assign T676 = $signed(30'h2769a939) * $signed(16'h0);
  assign T677 = T675[6'h2d:6'h2d];
  assign twiddle3_2_39_imag = T680 + T678;
  assign T678 = $signed(T679) / $signed(22'h100000);
  assign T679 = $signed(31'h39bd1c70) * $signed(16'hffff);
  assign T680 = {T683, T681};
  assign T681 = $signed(T682) / $signed(22'h100000);
  assign T682 = $signed(30'h24642bb3) * $signed(16'h0);
  assign T683 = T681[6'h2d:6'h2d];
  assign T684 = T383[1'h0:1'h0];
  assign T685 = T383[1'h1:1'h1];
  assign T686 = T383[2'h2:2'h2];
  assign T687 = T734 ? T712 : T688;
  assign T688 = T711 ? T701 : T689;
  assign T689 = T700 ? twiddle3_2_41_imag : twiddle3_2_40_imag;
  assign twiddle3_2_40_imag = T692 + T690;
  assign T690 = $signed(T691) / $signed(22'h100000);
  assign T691 = $signed(31'h383c0315) * $signed(16'hffff);
  assign T692 = {T695, T693};
  assign T693 = $signed(T694) / $signed(22'h100000);
  assign T694 = $signed(30'h217193da) * $signed(16'h0);
  assign T695 = T693[6'h2d:6'h2d];
  assign twiddle3_2_41_imag = T698 + T696;
  assign T696 = $signed(T697) / $signed(22'h100000);
  assign T697 = $signed(31'h36946c2f) * $signed(16'hffff);
  assign T698 = $signed(T699) / $signed(22'h100000);
  assign T699 = $signed(31'h5e93e62b) * $signed(16'h0);
  assign T700 = T383[1'h0:1'h0];
  assign T701 = T710 ? twiddle3_2_43_imag : twiddle3_2_42_imag;
  assign twiddle3_2_42_imag = T704 + T702;
  assign T702 = $signed(T703) / $signed(22'h100000);
  assign T703 = $signed(31'h34c779ab) * $signed(16'hffff);
  assign T704 = $signed(T705) / $signed(22'h100000);
  assign T705 = $signed(31'h5bcd18d2) * $signed(16'h0);
  assign twiddle3_2_43_imag = T708 + T706;
  assign T706 = $signed(T707) / $signed(22'h100000);
  assign T707 = $signed(31'h32d6670a) * $signed(16'hffff);
  assign T708 = $signed(T709) / $signed(22'h100000);
  assign T709 = $signed(31'h591f1255) * $signed(16'h0);
  assign T710 = T383[1'h0:1'h0];
  assign T711 = T383[1'h1:1'h1];
  assign T712 = T733 ? T723 : T713;
  assign T713 = T722 ? twiddle3_2_45_imag : twiddle3_2_44_imag;
  assign twiddle3_2_44_imag = T716 + T714;
  assign T714 = $signed(T715) / $signed(22'h100000);
  assign T715 = $signed(31'h30c28886) * $signed(16'hffff);
  assign T716 = $signed(T717) / $signed(22'h100000);
  assign T717 = $signed(31'h568ba843) * $signed(16'h0);
  assign twiddle3_2_45_imag = T720 + T718;
  assign T718 = $signed(T719) / $signed(22'h100000);
  assign T719 = $signed(31'h2e8d4a2c) * $signed(16'hffff);
  assign T720 = $signed(T721) / $signed(22'h100000);
  assign T721 = $signed(31'h54149df5) * $signed(16'h0);
  assign T722 = T383[1'h0:1'h0];
  assign T723 = T732 ? twiddle3_2_47_imag : twiddle3_2_46_imag;
  assign twiddle3_2_46_imag = T726 + T724;
  assign T724 = $signed(T725) / $signed(22'h100000);
  assign T725 = $signed(31'h2c382ede) * $signed(16'hffff);
  assign T726 = $signed(T727) / $signed(22'h100000);
  assign T727 = $signed(31'h51bba355) * $signed(16'h0);
  assign twiddle3_2_47_imag = T730 + T728;
  assign T728 = $signed(T729) / $signed(22'h100000);
  assign T729 = $signed(31'h29c4cf50) * $signed(16'hffff);
  assign T730 = $signed(T731) / $signed(22'h100000);
  assign T731 = $signed(31'h4f8253bf) * $signed(16'h0);
  assign T732 = T383[1'h0:1'h0];
  assign T733 = T383[1'h1:1'h1];
  assign T734 = T383[2'h2:2'h2];
  assign T735 = T383[2'h3:2'h3];
  assign T736 = T863 ? T793 : T737;
  assign T737 = T792 ? T762 : T738;
  assign T738 = T761 ? T749 : T739;
  assign T739 = T748 ? twiddle3_2_49_imag : twiddle3_2_48_imag;
  assign twiddle3_2_48_imag = T742 + T740;
  assign T740 = $signed(T741) / $signed(22'h100000);
  assign T741 = $signed(31'h2734d8ea) * $signed(16'hffff);
  assign T742 = $signed(T743) / $signed(22'h100000);
  assign T743 = $signed(31'h4d6a34de) * $signed(16'h0);
  assign twiddle3_2_49_imag = T746 + T744;
  assign T744 = $signed(T745) / $signed(22'h100000);
  assign T745 = $signed(31'h248a0caa) * $signed(16'hffff);
  assign T746 = $signed(T747) / $signed(22'h100000);
  assign T747 = $signed(31'h4b74b5a6) * $signed(16'h0);
  assign T748 = T383[1'h0:1'h0];
  assign T749 = T760 ? twiddle3_2_51_imag : twiddle3_2_50_imag;
  assign twiddle3_2_50_imag = T752 + T750;
  assign T750 = $signed(T751) / $signed(22'h100000);
  assign T751 = $signed(31'h21c63de7) * $signed(16'hffff);
  assign T752 = $signed(T753) / $signed(22'h100000);
  assign T753 = $signed(31'h49a32d5a) * $signed(16'h0);
  assign twiddle3_2_51_imag = T758 + T754;
  assign T754 = {T757, T755};
  assign T755 = $signed(T756) / $signed(22'h100000);
  assign T756 = $signed(30'h1eeb511b) * $signed(16'hffff);
  assign T757 = T755[6'h2d:6'h2d];
  assign T758 = $signed(T759) / $signed(22'h100000);
  assign T759 = $signed(31'h47f6da9c) * $signed(16'h0);
  assign T760 = T383[1'h0:1'h0];
  assign T761 = T383[1'h1:1'h1];
  assign T762 = T791 ? T777 : T763;
  assign T763 = T776 ? twiddle3_2_53_imag : twiddle3_2_52_imag;
  assign twiddle3_2_52_imag = T768 + T764;
  assign T764 = {T767, T765};
  assign T765 = $signed(T766) / $signed(22'h100000);
  assign T766 = $signed(30'h1bfb3a90) * $signed(16'hffff);
  assign T767 = T765[6'h2d:6'h2d];
  assign T768 = $signed(T769) / $signed(22'h100000);
  assign T769 = $signed(31'h4670e29a) * $signed(16'h0);
  assign twiddle3_2_53_imag = T774 + T770;
  assign T770 = {T773, T771};
  assign T771 = $signed(T772) / $signed(22'h100000);
  assign T772 = $signed(30'h18f7fd0d) * $signed(16'hffff);
  assign T773 = T771[6'h2d:6'h2d];
  assign T774 = $signed(T775) / $signed(22'h100000);
  assign T775 = $signed(31'h4512503e) * $signed(16'h0);
  assign T776 = T383[1'h0:1'h0];
  assign T777 = T790 ? twiddle3_2_55_imag : twiddle3_2_54_imag;
  assign twiddle3_2_54_imag = T782 + T778;
  assign T778 = {T781, T779};
  assign T779 = $signed(T780) / $signed(22'h100000);
  assign T780 = $signed(30'h15e3a874) * $signed(16'hffff);
  assign T781 = T779[6'h2d:6'h2d];
  assign T782 = $signed(T783) / $signed(22'h100000);
  assign T783 = $signed(31'h43dc137c) * $signed(16'h0);
  assign twiddle3_2_55_imag = T788 + T784;
  assign T784 = {T787, T785};
  assign T785 = $signed(T786) / $signed(22'h100000);
  assign T786 = $signed(30'h12c0585b) * $signed(16'hffff);
  assign T787 = T785[6'h2d:6'h2d];
  assign T788 = $signed(T789) / $signed(22'h100000);
  assign T789 = $signed(31'h42cf00ad) * $signed(16'h0);
  assign T790 = T383[1'h0:1'h0];
  assign T791 = T383[1'h1:1'h1];
  assign T792 = T383[2'h2:2'h2];
  assign T793 = T862 ? T828 : T794;
  assign T794 = T827 ? T811 : T795;
  assign T795 = T810 ? twiddle3_2_57_imag : twiddle3_2_56_imag;
  assign twiddle3_2_56_imag = T801 + T796;
  assign T796 = {T799, T797};
  assign T797 = $signed(T798) / $signed(22'h100000);
  assign T798 = $signed(29'hf903299) * $signed(16'hffff);
  assign T799 = T800 ? 2'h3 : 2'h0;
  assign T800 = T797[6'h2c:6'h2c];
  assign T801 = $signed(T802) / $signed(22'h100000);
  assign T802 = $signed(31'h41ebcffd) * $signed(16'h0);
  assign twiddle3_2_57_imag = T808 + T803;
  assign T803 = {T806, T804};
  assign T804 = $signed(T805) / $signed(22'h100000);
  assign T805 = $signed(29'hc5565ce) * $signed(16'hffff);
  assign T806 = T807 ? 2'h3 : 2'h0;
  assign T807 = T804[6'h2c:6'h2c];
  assign T808 = $signed(T809) / $signed(22'h100000);
  assign T809 = $signed(31'h41331ced) * $signed(16'h0);
  assign T810 = T383[1'h0:1'h0];
  assign T811 = T826 ? twiddle3_2_59_imag : twiddle3_2_58_imag;
  assign twiddle3_2_58_imag = T817 + T812;
  assign T812 = {T815, T813};
  assign T813 = $signed(T814) / $signed(22'h100000);
  assign T814 = $signed(29'h91227e2) * $signed(16'hffff);
  assign T815 = T816 ? 2'h3 : 2'h0;
  assign T816 = T813[6'h2c:6'h2c];
  assign T817 = $signed(T818) / $signed(22'h100000);
  assign T818 = $signed(31'h40a565e9) * $signed(16'h0);
  assign twiddle3_2_59_imag = T824 + T819;
  assign T819 = {T822, T820};
  assign T820 = $signed(T821) / $signed(22'h100000);
  assign T821 = $signed(28'h5c8b488) * $signed(16'hffff);
  assign T822 = T823 ? 3'h7 : 3'h0;
  assign T823 = T820[6'h2b:6'h2b];
  assign T824 = $signed(T825) / $signed(22'h100000);
  assign T825 = $signed(31'h40430bef) * $signed(16'h0);
  assign T826 = T383[1'h0:1'h0];
  assign T827 = T383[1'h1:1'h1];
  assign T828 = T861 ? T845 : T829;
  assign T829 = T844 ? twiddle3_2_61_imag : twiddle3_2_60_imag;
  assign twiddle3_2_60_imag = T835 + T830;
  assign T830 = {T833, T831};
  assign T831 = $signed(T832) / $signed(22'h100000);
  assign T832 = $signed(27'h27b4bb1) * $signed(16'hffff);
  assign T833 = T834 ? 4'hf : 4'h0;
  assign T834 = T831[6'h2a:6'h2a];
  assign T835 = $signed(T836) / $signed(22'h100000);
  assign T836 = $signed(31'h400c5251) * $signed(16'h0);
  assign twiddle3_2_61_imag = T842 + T837;
  assign T837 = {T840, T838};
  assign T838 = $signed(T839) / $signed(22'h100000);
  assign T839 = $signed(25'h12c3005) * $signed(16'hffff);
  assign T840 = T841 ? 6'h3f : 6'h0;
  assign T841 = T838[6'h28:6'h28];
  assign T842 = $signed(T843) / $signed(22'h100000);
  assign T843 = $signed(31'h40015e85) * $signed(16'h0);
  assign T844 = T383[1'h0:1'h0];
  assign T845 = T860 ? twiddle3_2_63_imag : twiddle3_2_62_imag;
  assign twiddle3_2_62_imag = T851 + T846;
  assign T846 = {T849, T847};
  assign T847 = $signed(T848) / $signed(22'h100000);
  assign T848 = $signed(28'hbdda552) * $signed(16'hffff);
  assign T849 = T850 ? 3'h7 : 3'h0;
  assign T850 = T847[6'h2b:6'h2b];
  assign T851 = $signed(T852) / $signed(22'h100000);
  assign T852 = $signed(31'h4022380a) * $signed(16'h0);
  assign twiddle3_2_63_imag = T858 + T853;
  assign T853 = {T856, T854};
  assign T854 = $signed(T855) / $signed(22'h100000);
  assign T855 = $signed(28'h891ef07) * $signed(16'hffff);
  assign T856 = T857 ? 3'h7 : 3'h0;
  assign T857 = T854[6'h2b:6'h2b];
  assign T858 = $signed(T859) / $signed(22'h100000);
  assign T859 = $signed(31'h406ec863) * $signed(16'h0);
  assign T860 = T383[1'h0:1'h0];
  assign T861 = T383[1'h1:1'h1];
  assign T862 = T383[2'h2:2'h2];
  assign T863 = T383[2'h3:2'h3];
  assign T864 = T383[3'h4:3'h4];
  assign T865 = T619[6'h2e:6'h2e];
  assign T866 = T383[3'h5:3'h5];
  assign T867 = {T984, T868};
  assign T868 = T983 ? twiddle3_2_80_imag : T869;
  assign T869 = T978 ? T932 : T870;
  assign T870 = T931 ? T903 : T871;
  assign T871 = T902 ? T888 : T872;
  assign T872 = T887 ? twiddle3_2_65_imag : twiddle3_2_64_imag;
  assign twiddle3_2_64_imag = T878 + T873;
  assign T873 = {T876, T874};
  assign T874 = $signed(T875) / $signed(22'h100000);
  assign T875 = $signed(29'h154b4ea1) * $signed(16'hffff);
  assign T876 = T877 ? 2'h3 : 2'h0;
  assign T877 = T874[6'h2c:6'h2c];
  assign T878 = $signed(T879) / $signed(22'h100000);
  assign T879 = $signed(31'h40e6db28) * $signed(16'h0);
  assign twiddle3_2_65_imag = T885 + T880;
  assign T880 = {T883, T881};
  assign T881 = $signed(T882) / $signed(22'h100000);
  assign T882 = $signed(29'h120c0223) * $signed(16'hffff);
  assign T883 = T884 ? 2'h3 : 2'h0;
  assign T884 = T881[6'h2c:6'h2c];
  assign T885 = $signed(T886) / $signed(22'h100000);
  assign T886 = $signed(31'h418a1e2b) * $signed(16'h0);
  assign T887 = T383[1'h0:1'h0];
  assign T888 = T901 ? twiddle3_2_67_imag : twiddle3_2_66_imag;
  assign twiddle3_2_66_imag = T893 + T889;
  assign T889 = {T892, T890};
  assign T890 = $signed(T891) / $signed(22'h100000);
  assign T891 = $signed(30'h2ed6428a) * $signed(16'hffff);
  assign T892 = T890[6'h2d:6'h2d];
  assign T893 = $signed(T894) / $signed(22'h100000);
  assign T894 = $signed(31'h425821ac) * $signed(16'h0);
  assign twiddle3_2_67_imag = T899 + T895;
  assign T895 = {T898, T896};
  assign T896 = $signed(T897) / $signed(22'h100000);
  assign T897 = $signed(30'h2bac424d) * $signed(16'hffff);
  assign T898 = T896[6'h2d:6'h2d];
  assign T899 = $signed(T900) / $signed(22'h100000);
  assign T900 = $signed(31'h435058a9) * $signed(16'h0);
  assign T901 = T383[1'h0:1'h0];
  assign T902 = T383[1'h1:1'h1];
  assign T903 = T930 ? T918 : T904;
  assign T904 = T917 ? twiddle3_2_69_imag : twiddle3_2_68_imag;
  assign twiddle3_2_68_imag = T909 + T905;
  assign T905 = {T908, T906};
  assign T906 = $signed(T907) / $signed(22'h100000);
  assign T907 = $signed(30'h28902bd4) * $signed(16'hffff);
  assign T908 = T906[6'h2d:6'h2d];
  assign T909 = $signed(T910) / $signed(22'h100000);
  assign T910 = $signed(31'h4472193c) * $signed(16'h0);
  assign twiddle3_2_69_imag = T915 + T911;
  assign T911 = {T914, T912};
  assign T912 = $signed(T913) / $signed(22'h100000);
  assign T913 = $signed(30'h25842006) * $signed(16'hffff);
  assign T914 = T912[6'h2d:6'h2d];
  assign T915 = $signed(T916) / $signed(22'h100000);
  assign T916 = $signed(31'h45bc9d14) * $signed(16'h0);
  assign T917 = T383[1'h0:1'h0];
  assign T918 = T929 ? twiddle3_2_71_imag : twiddle3_2_70_imag;
  assign twiddle3_2_70_imag = T923 + T919;
  assign T919 = {T922, T920};
  assign T920 = $signed(T921) / $signed(22'h100000);
  assign T921 = $signed(30'h228a34cc) * $signed(16'hffff);
  assign T922 = T920[6'h2d:6'h2d];
  assign T923 = $signed(T924) / $signed(22'h100000);
  assign T924 = $signed(31'h472f01f5) * $signed(16'h0);
  assign twiddle3_2_71_imag = T927 + T925;
  assign T925 = $signed(T926) / $signed(22'h100000);
  assign T926 = $signed(31'h5fa473a7) * $signed(16'hffff);
  assign T927 = $signed(T928) / $signed(22'h100000);
  assign T928 = $signed(31'h48c84a5b) * $signed(16'h0);
  assign T929 = T383[1'h0:1'h0];
  assign T930 = T383[1'h1:1'h1];
  assign T931 = T383[2'h2:2'h2];
  assign T932 = T977 ? T955 : T933;
  assign T933 = T954 ? T944 : T934;
  assign T934 = T943 ? twiddle3_2_73_imag : twiddle3_2_72_imag;
  assign twiddle3_2_72_imag = T937 + T935;
  assign T935 = $signed(T936) / $signed(22'h100000);
  assign T936 = $signed(31'h5cd4d84c) * $signed(16'hffff);
  assign T937 = $signed(T938) / $signed(22'h100000);
  assign T938 = $signed(31'h4a875e22) * $signed(16'h0);
  assign twiddle3_2_73_imag = T941 + T939;
  assign T939 = $signed(T940) / $signed(22'h100000);
  assign T940 = $signed(31'h5a1d4f46) * $signed(16'hffff);
  assign T941 = $signed(T942) / $signed(22'h100000);
  assign T942 = $signed(31'h4c6b0b48) * $signed(16'h0);
  assign T943 = T383[1'h0:1'h0];
  assign T944 = T953 ? twiddle3_2_75_imag : twiddle3_2_74_imag;
  assign twiddle3_2_74_imag = T947 + T945;
  assign T945 = $signed(T946) / $signed(22'h100000);
  assign T946 = $signed(31'h577fb4a6) * $signed(16'hffff);
  assign T947 = $signed(T948) / $signed(22'h100000);
  assign T948 = $signed(31'h4e7206bd) * $signed(16'h0);
  assign twiddle3_2_75_imag = T951 + T949;
  assign T949 = $signed(T950) / $signed(22'h100000);
  assign T950 = $signed(31'h54fdd2bf) * $signed(16'hffff);
  assign T951 = $signed(T952) / $signed(22'h100000);
  assign T952 = $signed(31'h509aed49) * $signed(16'h0);
  assign T953 = T383[1'h0:1'h0];
  assign T954 = T383[1'h1:1'h1];
  assign T955 = T976 ? T966 : T956;
  assign T956 = T965 ? twiddle3_2_77_imag : twiddle3_2_76_imag;
  assign twiddle3_2_76_imag = T959 + T957;
  assign T957 = $signed(T958) / $signed(22'h100000);
  assign T958 = $signed(31'h529960e8) * $signed(16'hffff);
  assign T959 = $signed(T960) / $signed(22'h100000);
  assign T960 = $signed(31'h52e4447b) * $signed(16'h0);
  assign twiddle3_2_77_imag = T963 + T961;
  assign T961 = $signed(T962) / $signed(22'h100000);
  assign T962 = $signed(31'h50540254) * $signed(16'hffff);
  assign T963 = $signed(T964) / $signed(22'h100000);
  assign T964 = $signed(31'h554c7bad) * $signed(16'h0);
  assign T965 = T383[1'h0:1'h0];
  assign T966 = T975 ? twiddle3_2_79_imag : twiddle3_2_78_imag;
  assign twiddle3_2_78_imag = T969 + T967;
  assign T967 = $signed(T968) / $signed(22'h100000);
  assign T968 = $signed(31'h4e2f44f0) * $signed(16'hffff);
  assign T969 = $signed(T970) / $signed(22'h100000);
  assign T970 = $signed(31'h57d1ed19) * $signed(16'h0);
  assign twiddle3_2_79_imag = T973 + T971;
  assign T971 = $signed(T972) / $signed(22'h100000);
  assign T972 = $signed(31'h4c2ca054) * $signed(16'hffff);
  assign T973 = $signed(T974) / $signed(22'h100000);
  assign T974 = $signed(31'h5a72def6) * $signed(16'h0);
  assign T975 = T383[1'h0:1'h0];
  assign T976 = T383[1'h1:1'h1];
  assign T977 = T383[2'h2:2'h2];
  assign T978 = T383[2'h3:2'h3];
  assign twiddle3_2_80_imag = T981 + T979;
  assign T979 = $signed(T980) / $signed(22'h100000);
  assign T980 = $signed(31'h4a4d74c1) * $signed(16'hffff);
  assign T981 = $signed(T982) / $signed(22'h100000);
  assign T982 = $signed(31'h5d2d84aa) * $signed(16'h0);
  assign T983 = T383[3'h4:3'h4];
  assign T984 = T868[6'h2e:6'h2e];
  assign T985 = T383[3'h6:3'h6];
  assign io_t3_2out_real = T986;
  assign T986 = T987[4'hf:1'h0];
  assign T987 = T1611 ? T1493 : T988;
  assign T988 = T1492 ? T1244 : T989;
  assign T989 = T1243 ? T1119 : T990;
  assign T990 = T1118 ? T1064 : T991;
  assign T991 = T1063 ? T1030 : T992;
  assign T992 = T1029 ? T1011 : T993;
  assign T993 = T1010 ? T1001 : twiddle3_2_0_real;
  assign twiddle3_2_0_real = T999 + T994;
  assign T994 = {T997, T995};
  assign T995 = $signed(T996) / $signed(22'h100000);
  assign T996 = $signed(1'h0) * $signed(16'h0);
  assign T997 = T998 ? 31'h7fffffff : 31'h0;
  assign T998 = T995[5'h10:5'h10];
  assign T999 = $signed(T1000) / $signed(22'h100000);
  assign T1000 = $signed(32'h40000000) * $signed(16'h1);
  assign T1001 = {T1009, twiddle3_2_1_real};
  assign twiddle3_2_1_real = T1007 + T1002;
  assign T1002 = {T1005, T1003};
  assign T1003 = $signed(T1004) / $signed(22'h100000);
  assign T1004 = $signed(27'h34ee54e) * $signed(16'h0);
  assign T1005 = T1006 ? 4'hf : 4'h0;
  assign T1006 = T1003[6'h2a:6'h2a];
  assign T1007 = $signed(T1008) / $signed(22'h100000);
  assign T1008 = $signed(31'h3fea18df) * $signed(16'h1);
  assign T1009 = twiddle3_2_1_real[6'h2e:6'h2e];
  assign T1010 = T383[1'h0:1'h0];
  assign T1011 = {T1028, T1012};
  assign T1012 = T1027 ? twiddle3_2_3_real : twiddle3_2_2_real;
  assign twiddle3_2_2_real = T1018 + T1013;
  assign T1013 = {T1016, T1014};
  assign T1014 = $signed(T1015) / $signed(22'h100000);
  assign T1015 = $signed(28'h69b86f1) * $signed(16'h0);
  assign T1016 = T1017 ? 3'h7 : 3'h0;
  assign T1017 = T1014[6'h2b:6'h2b];
  assign T1018 = $signed(T1019) / $signed(22'h100000);
  assign T1019 = $signed(31'h3fa8727d) * $signed(16'h1);
  assign twiddle3_2_3_real = T1025 + T1020;
  assign T1020 = {T1023, T1021};
  assign T1021 = $signed(T1022) / $signed(22'h100000);
  assign T1022 = $signed(29'h9e3a2ca) * $signed(16'h0);
  assign T1023 = T1024 ? 2'h3 : 2'h0;
  assign T1024 = T1021[6'h2c:6'h2c];
  assign T1025 = $signed(T1026) / $signed(22'h100000);
  assign T1026 = $signed(31'h3f3b39c7) * $signed(16'h1);
  assign T1027 = T383[1'h0:1'h0];
  assign T1028 = T1012[6'h2e:6'h2e];
  assign T1029 = T383[1'h1:1'h1];
  assign T1030 = {T1062, T1031};
  assign T1031 = T1061 ? T1047 : T1032;
  assign T1032 = T1046 ? twiddle3_2_5_real : twiddle3_2_4_real;
  assign twiddle3_2_4_real = T1038 + T1033;
  assign T1033 = {T1036, T1034};
  assign T1034 = $signed(T1035) / $signed(22'h100000);
  assign T1035 = $signed(29'hd24f9d3) * $signed(16'h0);
  assign T1036 = T1037 ? 2'h3 : 2'h0;
  assign T1037 = T1034[6'h2c:6'h2c];
  assign T1038 = $signed(T1039) / $signed(22'h100000);
  assign T1039 = $signed(31'h3ea2b980) * $signed(16'h1);
  assign twiddle3_2_5_real = T1044 + T1040;
  assign T1040 = {T1043, T1041};
  assign T1041 = $signed(T1042) / $signed(22'h100000);
  assign T1042 = $signed(30'h105d51a8) * $signed(16'h0);
  assign T1043 = T1041[6'h2d:6'h2d];
  assign T1044 = $signed(T1045) / $signed(22'h100000);
  assign T1045 = $signed(31'h3ddf5a09) * $signed(16'h1);
  assign T1046 = T383[1'h0:1'h0];
  assign T1047 = T1060 ? twiddle3_2_7_real : twiddle3_2_6_real;
  assign twiddle3_2_6_real = T1052 + T1048;
  assign T1048 = {T1051, T1049};
  assign T1049 = $signed(T1050) / $signed(22'h100000);
  assign T1050 = $signed(30'h138a760d) * $signed(16'h0);
  assign T1051 = T1049[6'h2d:6'h2d];
  assign T1052 = $signed(T1053) / $signed(22'h100000);
  assign T1053 = $signed(31'h3cf1a11d) * $signed(16'h1);
  assign twiddle3_2_7_real = T1058 + T1054;
  assign T1054 = {T1057, T1055};
  assign T1055 = $signed(T1056) / $signed(22'h100000);
  assign T1056 = $signed(30'h16aa3a72) * $signed(16'h0);
  assign T1057 = T1055[6'h2d:6'h2d];
  assign T1058 = $signed(T1059) / $signed(22'h100000);
  assign T1059 = $signed(31'h3bda3171) * $signed(16'h1);
  assign T1060 = T383[1'h0:1'h0];
  assign T1061 = T383[1'h1:1'h1];
  assign T1062 = T1031[6'h2e:6'h2e];
  assign T1063 = T383[2'h2:2'h2];
  assign T1064 = {T1117, T1065};
  assign T1065 = T1116 ? T1094 : T1066;
  assign T1066 = T1093 ? T1081 : T1067;
  assign T1067 = T1080 ? twiddle3_2_9_real : twiddle3_2_8_real;
  assign twiddle3_2_8_real = T1072 + T1068;
  assign T1068 = {T1071, T1069};
  assign T1069 = $signed(T1070) / $signed(22'h100000);
  assign T1070 = $signed(30'h19ba7b6c) * $signed(16'h0);
  assign T1071 = T1069[6'h2d:6'h2d];
  assign T1072 = $signed(T1073) / $signed(22'h100000);
  assign T1073 = $signed(31'h3a99ca4a) * $signed(16'h1);
  assign twiddle3_2_9_real = T1078 + T1074;
  assign T1074 = {T1077, T1075};
  assign T1075 = $signed(T1076) / $signed(22'h100000);
  assign T1076 = $signed(30'h1cb92032) * $signed(16'h0);
  assign T1077 = T1075[6'h2d:6'h2d];
  assign T1078 = $signed(T1079) / $signed(22'h100000);
  assign T1079 = $signed(31'h393146f5) * $signed(16'h1);
  assign T1080 = T383[1'h0:1'h0];
  assign T1081 = T1092 ? twiddle3_2_11_real : twiddle3_2_10_real;
  assign twiddle3_2_10_real = T1086 + T1082;
  assign T1082 = {T1085, T1083};
  assign T1083 = $signed(T1084) / $signed(22'h100000);
  assign T1084 = $signed(30'h1fa41c05) * $signed(16'h0);
  assign T1085 = T1083[6'h2d:6'h2d];
  assign T1086 = $signed(T1087) / $signed(22'h100000);
  assign T1087 = $signed(31'h37a19e34) * $signed(16'h1);
  assign twiddle3_2_11_real = T1090 + T1088;
  assign T1088 = $signed(T1089) / $signed(22'h100000);
  assign T1089 = $signed(31'h22796f9d) * $signed(16'h0);
  assign T1090 = $signed(T1091) / $signed(22'h100000);
  assign T1091 = $signed(31'h35ebe194) * $signed(16'h1);
  assign T1092 = T383[1'h0:1'h0];
  assign T1093 = T383[1'h1:1'h1];
  assign T1094 = T1115 ? T1105 : T1095;
  assign T1095 = T1104 ? twiddle3_2_13_real : twiddle3_2_12_real;
  assign twiddle3_2_12_real = T1098 + T1096;
  assign T1096 = $signed(T1097) / $signed(22'h100000);
  assign T1097 = $signed(31'h25372a85) * $signed(16'h0);
  assign T1098 = $signed(T1099) / $signed(22'h100000);
  assign T1099 = $signed(31'h34113cb3) * $signed(16'h1);
  assign twiddle3_2_13_real = T1102 + T1100;
  assign T1100 = $signed(T1101) / $signed(22'h100000);
  assign T1101 = $signed(31'h27db6c6d) * $signed(16'h0);
  assign T1102 = $signed(T1103) / $signed(22'h100000);
  assign T1103 = $signed(31'h3212f472) * $signed(16'h1);
  assign T1104 = T383[1'h0:1'h0];
  assign T1105 = T1114 ? twiddle3_2_15_real : twiddle3_2_14_real;
  assign twiddle3_2_14_real = T1108 + T1106;
  assign T1106 = $signed(T1107) / $signed(22'h100000);
  assign T1107 = $signed(31'h2a646676) * $signed(16'h0);
  assign T1108 = $signed(T1109) / $signed(22'h100000);
  assign T1109 = $signed(31'h2ff26615) * $signed(16'h1);
  assign twiddle3_2_15_real = T1112 + T1110;
  assign T1110 = $signed(T1111) / $signed(22'h100000);
  assign T1111 = $signed(31'h2cd05c6c) * $signed(16'h0);
  assign T1112 = $signed(T1113) / $signed(22'h100000);
  assign T1113 = $signed(31'h2db10657) * $signed(16'h1);
  assign T1114 = T383[1'h0:1'h0];
  assign T1115 = T383[1'h1:1'h1];
  assign T1116 = T383[2'h2:2'h2];
  assign T1117 = T1065[6'h2e:6'h2e];
  assign T1118 = T383[2'h3:2'h3];
  assign T1119 = {T1242, T1120};
  assign T1120 = T1241 ? T1173 : T1121;
  assign T1121 = T1172 ? T1144 : T1122;
  assign T1122 = T1143 ? T1133 : T1123;
  assign T1123 = T1132 ? twiddle3_2_17_real : twiddle3_2_16_real;
  assign twiddle3_2_16_real = T1126 + T1124;
  assign T1124 = $signed(T1125) / $signed(22'h100000);
  assign T1125 = $signed(31'h2f1da5f8) * $signed(16'h0);
  assign T1126 = $signed(T1127) / $signed(22'h100000);
  assign T1127 = $signed(31'h2b506069) * $signed(16'h1);
  assign twiddle3_2_17_real = T1130 + T1128;
  assign T1128 = $signed(T1129) / $signed(22'h100000);
  assign T1129 = $signed(31'h314aafc2) * $signed(16'h0);
  assign T1130 = $signed(T1131) / $signed(22'h100000);
  assign T1131 = $signed(31'h28d214e4) * $signed(16'h1);
  assign T1132 = T383[1'h0:1'h0];
  assign T1133 = T1142 ? twiddle3_2_19_real : twiddle3_2_18_real;
  assign twiddle3_2_18_real = T1136 + T1134;
  assign T1134 = $signed(T1135) / $signed(22'h100000);
  assign T1135 = $signed(31'h3355fc84) * $signed(16'h0);
  assign T1136 = $signed(T1137) / $signed(22'h100000);
  assign T1137 = $signed(31'h2637d8ab) * $signed(16'h1);
  assign twiddle3_2_19_real = T1140 + T1138;
  assign T1138 = $signed(T1139) / $signed(22'h100000);
  assign T1139 = $signed(31'h353e260f) * $signed(16'h0);
  assign T1140 = $signed(T1141) / $signed(22'h100000);
  assign T1141 = $signed(31'h238373c3) * $signed(16'h1);
  assign T1142 = T383[1'h0:1'h0];
  assign T1143 = T383[1'h1:1'h1];
  assign T1144 = T1171 ? T1157 : T1145;
  assign T1145 = T1156 ? twiddle3_2_21_real : twiddle3_2_20_real;
  assign twiddle3_2_20_real = T1148 + T1146;
  assign T1146 = $signed(T1147) / $signed(22'h100000);
  assign T1147 = $signed(31'h3701de44) * $signed(16'h0);
  assign T1148 = $signed(T1149) / $signed(22'h100000);
  assign T1149 = $signed(31'h20b6c016) * $signed(16'h1);
  assign twiddle3_2_21_real = T1152 + T1150;
  assign T1150 = $signed(T1151) / $signed(22'h100000);
  assign T1151 = $signed(31'h389feff1) * $signed(16'h0);
  assign T1152 = {T1155, T1153};
  assign T1153 = $signed(T1154) / $signed(22'h100000);
  assign T1154 = $signed(30'h1dd3a832) * $signed(16'h1);
  assign T1155 = T1153[6'h2d:6'h2d];
  assign T1156 = T383[1'h0:1'h0];
  assign T1157 = T1170 ? twiddle3_2_23_real : twiddle3_2_22_real;
  assign twiddle3_2_22_real = T1160 + T1158;
  assign T1158 = $signed(T1159) / $signed(22'h100000);
  assign T1159 = $signed(31'h3a173fae) * $signed(16'h0);
  assign T1160 = {T1163, T1161};
  assign T1161 = $signed(T1162) / $signed(22'h100000);
  assign T1162 = $signed(30'h1adc25fb) * $signed(16'h1);
  assign T1163 = T1161[6'h2d:6'h2d];
  assign twiddle3_2_23_real = T1166 + T1164;
  assign T1164 = $signed(T1165) / $signed(22'h100000);
  assign T1165 = $signed(31'h3b66cc97) * $signed(16'h0);
  assign T1166 = {T1169, T1167};
  assign T1167 = $signed(T1168) / $signed(22'h100000);
  assign T1168 = $signed(30'h17d2414a) * $signed(16'h1);
  assign T1169 = T1167[6'h2d:6'h2d];
  assign T1170 = T383[1'h0:1'h0];
  assign T1171 = T383[1'h1:1'h1];
  assign T1172 = T383[2'h2:2'h2];
  assign T1173 = T1240 ? T1206 : T1174;
  assign T1174 = T1205 ? T1189 : T1175;
  assign T1175 = T1188 ? twiddle3_2_25_real : twiddle3_2_24_real;
  assign twiddle3_2_24_real = T1178 + T1176;
  assign T1176 = $signed(T1177) / $signed(22'h100000);
  assign T1177 = $signed(31'h3c8db0ff) * $signed(16'h0);
  assign T1178 = {T1181, T1179};
  assign T1179 = $signed(T1180) / $signed(22'h100000);
  assign T1180 = $signed(30'h14b80e91) * $signed(16'h1);
  assign T1181 = T1179[6'h2d:6'h2d];
  assign twiddle3_2_25_real = T1184 + T1182;
  assign T1182 = $signed(T1183) / $signed(22'h100000);
  assign T1183 = $signed(31'h3d8b2310) * $signed(16'h0);
  assign T1184 = {T1187, T1185};
  assign T1185 = $signed(T1186) / $signed(22'h100000);
  assign T1186 = $signed(30'h118fad69) * $signed(16'h1);
  assign T1187 = T1185[6'h2d:6'h2d];
  assign T1188 = T383[1'h0:1'h0];
  assign T1189 = T1204 ? twiddle3_2_27_real : twiddle3_2_26_real;
  assign twiddle3_2_26_real = T1192 + T1190;
  assign T1190 = $signed(T1191) / $signed(22'h100000);
  assign T1191 = $signed(31'h3e5e754f) * $signed(16'h0);
  assign T1192 = {T1195, T1193};
  assign T1193 = $signed(T1194) / $signed(22'h100000);
  assign T1194 = $signed(29'he5b4720) * $signed(16'h1);
  assign T1195 = T1196 ? 2'h3 : 2'h0;
  assign T1196 = T1193[6'h2c:6'h2c];
  assign twiddle3_2_27_real = T1199 + T1197;
  assign T1197 = $signed(T1198) / $signed(22'h100000);
  assign T1198 = $signed(31'h3f071719) * $signed(16'h0);
  assign T1199 = {T1202, T1200};
  assign T1200 = $signed(T1201) / $signed(22'h100000);
  assign T1201 = $signed(29'hb1d0d3f) * $signed(16'h1);
  assign T1202 = T1203 ? 2'h3 : 2'h0;
  assign T1203 = T1200[6'h2c:6'h2c];
  assign T1204 = T383[1'h0:1'h0];
  assign T1205 = T383[1'h1:1'h1];
  assign T1206 = T1239 ? T1223 : T1207;
  assign T1207 = T1222 ? twiddle3_2_29_real : twiddle3_2_28_real;
  assign twiddle3_2_28_real = T1210 + T1208;
  assign T1208 = $signed(T1209) / $signed(22'h100000);
  assign T1209 = $signed(31'h3f849500) * $signed(16'h0);
  assign T1210 = {T1213, T1211};
  assign T1211 = $signed(T1212) / $signed(22'h100000);
  assign T1212 = $signed(28'h7d73808) * $signed(16'h1);
  assign T1213 = T1214 ? 3'h7 : 3'h0;
  assign T1214 = T1211[6'h2b:6'h2b];
  assign twiddle3_2_29_real = T1217 + T1215;
  assign T1215 = $signed(T1216) / $signed(22'h100000);
  assign T1216 = $signed(31'h3fd69921) * $signed(16'h0);
  assign T1217 = {T1220, T1218};
  assign T1218 = $signed(T1219) / $signed(22'h100000);
  assign T1219 = $signed(28'h48c04f3) * $signed(16'h1);
  assign T1220 = T1221 ? 3'h7 : 3'h0;
  assign T1221 = T1218[6'h2b:6'h2b];
  assign T1222 = T383[1'h0:1'h0];
  assign T1223 = T1238 ? twiddle3_2_31_real : twiddle3_2_30_real;
  assign twiddle3_2_30_real = T1226 + T1224;
  assign T1224 = $signed(T1225) / $signed(22'h100000);
  assign T1225 = $signed(31'h3ffceb58) * $signed(16'h0);
  assign T1226 = {T1229, T1227};
  assign T1227 = $signed(T1228) / $signed(22'h100000);
  assign T1228 = $signed(26'h13db523) * $signed(16'h1);
  assign T1229 = T1230 ? 5'h1f : 5'h0;
  assign T1230 = T1227[6'h29:6'h29];
  assign twiddle3_2_31_real = T1233 + T1231;
  assign T1231 = $signed(T1232) / $signed(22'h100000);
  assign T1232 = $signed(31'h3ff7716b) * $signed(16'h0);
  assign T1233 = {T1236, T1234};
  assign T1234 = $signed(T1235) / $signed(22'h100000);
  assign T1235 = $signed(27'h5ee8bdf) * $signed(16'h1);
  assign T1236 = T1237 ? 4'hf : 4'h0;
  assign T1237 = T1234[6'h2a:6'h2a];
  assign T1238 = T383[1'h0:1'h0];
  assign T1239 = T383[1'h1:1'h1];
  assign T1240 = T383[2'h2:2'h2];
  assign T1241 = T383[2'h3:2'h3];
  assign T1242 = T1120[6'h2e:6'h2e];
  assign T1243 = T383[3'h4:3'h4];
  assign T1244 = {T1491, T1245};
  assign T1245 = T1490 ? T1362 : T1246;
  assign T1246 = T1361 ? T1313 : T1247;
  assign T1247 = T1312 ? T1282 : T1248;
  assign T1248 = T1281 ? T1265 : T1249;
  assign T1249 = T1264 ? twiddle3_2_33_real : twiddle3_2_32_real;
  assign twiddle3_2_32_real = T1252 + T1250;
  assign T1250 = $signed(T1251) / $signed(22'h100000);
  assign T1251 = $signed(31'h3fc62f18) * $signed(16'h0);
  assign T1252 = {T1255, T1253};
  assign T1253 = $signed(T1254) / $signed(22'h100000);
  assign T1254 = $signed(28'haa0ccff) * $signed(16'h1);
  assign T1255 = T1256 ? 3'h7 : 3'h0;
  assign T1256 = T1253[6'h2b:6'h2b];
  assign twiddle3_2_33_real = T1259 + T1257;
  assign T1257 = $signed(T1258) / $signed(22'h100000);
  assign T1258 = $signed(31'h3f694618) * $signed(16'h0);
  assign T1259 = {T1262, T1260};
  assign T1260 = $signed(T1261) / $signed(22'h100000);
  assign T1261 = $signed(29'h1756bb64) * $signed(16'h1);
  assign T1262 = T1263 ? 2'h3 : 2'h0;
  assign T1263 = T1260[6'h2c:6'h2c];
  assign T1264 = T383[1'h0:1'h0];
  assign T1265 = T1280 ? twiddle3_2_35_real : twiddle3_2_34_real;
  assign twiddle3_2_34_real = T1268 + T1266;
  assign T1266 = $signed(T1267) / $signed(22'h100000);
  assign T1267 = $signed(31'h3ee0f602) * $signed(16'h0);
  assign T1268 = {T1271, T1269};
  assign T1269 = $signed(T1270) / $signed(22'h100000);
  assign T1270 = $signed(29'h1412976d) * $signed(16'h1);
  assign T1271 = T1272 ? 2'h3 : 2'h0;
  assign T1272 = T1269[6'h2c:6'h2c];
  assign twiddle3_2_35_real = T1275 + T1273;
  assign T1273 = $signed(T1274) / $signed(22'h100000);
  assign T1274 = $signed(31'h3e2d9c23) * $signed(16'h0);
  assign T1275 = {T1278, T1276};
  assign T1276 = $signed(T1277) / $signed(22'h100000);
  assign T1277 = $signed(29'h10d69d68) * $signed(16'h1);
  assign T1278 = T1279 ? 2'h3 : 2'h0;
  assign T1279 = T1276[6'h2c:6'h2c];
  assign T1280 = T383[1'h0:1'h0];
  assign T1281 = T383[1'h1:1'h1];
  assign T1282 = T1311 ? T1297 : T1283;
  assign T1283 = T1296 ? twiddle3_2_37_real : twiddle3_2_36_real;
  assign twiddle3_2_36_real = T1286 + T1284;
  assign T1284 = $signed(T1285) / $signed(22'h100000);
  assign T1285 = $signed(31'h3d4fb33e) * $signed(16'h0);
  assign T1286 = {T1289, T1287};
  assign T1287 = $signed(T1288) / $signed(22'h100000);
  assign T1288 = $signed(30'h2da5040e) * $signed(16'h1);
  assign T1289 = T1287[6'h2d:6'h2d];
  assign twiddle3_2_37_real = T1292 + T1290;
  assign T1290 = $signed(T1291) / $signed(22'h100000);
  assign T1291 = $signed(31'h3c47d336) * $signed(16'h0);
  assign T1292 = {T1295, T1293};
  assign T1293 = $signed(T1294) / $signed(22'h100000);
  assign T1294 = $signed(30'h2a7ffafd) * $signed(16'h1);
  assign T1295 = T1293[6'h2d:6'h2d];
  assign T1296 = T383[1'h0:1'h0];
  assign T1297 = T1310 ? twiddle3_2_39_real : twiddle3_2_38_real;
  assign twiddle3_2_38_real = T1300 + T1298;
  assign T1298 = $signed(T1299) / $signed(22'h100000);
  assign T1299 = $signed(31'h3b16b0a8) * $signed(16'h0);
  assign T1300 = {T1303, T1301};
  assign T1301 = $signed(T1302) / $signed(22'h100000);
  assign T1302 = $signed(30'h2769a939) * $signed(16'h1);
  assign T1303 = T1301[6'h2d:6'h2d];
  assign twiddle3_2_39_real = T1306 + T1304;
  assign T1304 = $signed(T1305) / $signed(22'h100000);
  assign T1305 = $signed(31'h39bd1c70) * $signed(16'h0);
  assign T1306 = {T1309, T1307};
  assign T1307 = $signed(T1308) / $signed(22'h100000);
  assign T1308 = $signed(30'h24642bb3) * $signed(16'h1);
  assign T1309 = T1307[6'h2d:6'h2d];
  assign T1310 = T383[1'h0:1'h0];
  assign T1311 = T383[1'h1:1'h1];
  assign T1312 = T383[2'h2:2'h2];
  assign T1313 = T1360 ? T1338 : T1314;
  assign T1314 = T1337 ? T1327 : T1315;
  assign T1315 = T1326 ? twiddle3_2_41_real : twiddle3_2_40_real;
  assign twiddle3_2_40_real = T1318 + T1316;
  assign T1316 = $signed(T1317) / $signed(22'h100000);
  assign T1317 = $signed(31'h383c0315) * $signed(16'h0);
  assign T1318 = {T1321, T1319};
  assign T1319 = $signed(T1320) / $signed(22'h100000);
  assign T1320 = $signed(30'h217193da) * $signed(16'h1);
  assign T1321 = T1319[6'h2d:6'h2d];
  assign twiddle3_2_41_real = T1324 + T1322;
  assign T1322 = $signed(T1323) / $signed(22'h100000);
  assign T1323 = $signed(31'h36946c2f) * $signed(16'h0);
  assign T1324 = $signed(T1325) / $signed(22'h100000);
  assign T1325 = $signed(31'h5e93e62b) * $signed(16'h1);
  assign T1326 = T383[1'h0:1'h0];
  assign T1327 = T1336 ? twiddle3_2_43_real : twiddle3_2_42_real;
  assign twiddle3_2_42_real = T1330 + T1328;
  assign T1328 = $signed(T1329) / $signed(22'h100000);
  assign T1329 = $signed(31'h34c779ab) * $signed(16'h0);
  assign T1330 = $signed(T1331) / $signed(22'h100000);
  assign T1331 = $signed(31'h5bcd18d2) * $signed(16'h1);
  assign twiddle3_2_43_real = T1334 + T1332;
  assign T1332 = $signed(T1333) / $signed(22'h100000);
  assign T1333 = $signed(31'h32d6670a) * $signed(16'h0);
  assign T1334 = $signed(T1335) / $signed(22'h100000);
  assign T1335 = $signed(31'h591f1255) * $signed(16'h1);
  assign T1336 = T383[1'h0:1'h0];
  assign T1337 = T383[1'h1:1'h1];
  assign T1338 = T1359 ? T1349 : T1339;
  assign T1339 = T1348 ? twiddle3_2_45_real : twiddle3_2_44_real;
  assign twiddle3_2_44_real = T1342 + T1340;
  assign T1340 = $signed(T1341) / $signed(22'h100000);
  assign T1341 = $signed(31'h30c28886) * $signed(16'h0);
  assign T1342 = $signed(T1343) / $signed(22'h100000);
  assign T1343 = $signed(31'h568ba843) * $signed(16'h1);
  assign twiddle3_2_45_real = T1346 + T1344;
  assign T1344 = $signed(T1345) / $signed(22'h100000);
  assign T1345 = $signed(31'h2e8d4a2c) * $signed(16'h0);
  assign T1346 = $signed(T1347) / $signed(22'h100000);
  assign T1347 = $signed(31'h54149df5) * $signed(16'h1);
  assign T1348 = T383[1'h0:1'h0];
  assign T1349 = T1358 ? twiddle3_2_47_real : twiddle3_2_46_real;
  assign twiddle3_2_46_real = T1352 + T1350;
  assign T1350 = $signed(T1351) / $signed(22'h100000);
  assign T1351 = $signed(31'h2c382ede) * $signed(16'h0);
  assign T1352 = $signed(T1353) / $signed(22'h100000);
  assign T1353 = $signed(31'h51bba355) * $signed(16'h1);
  assign twiddle3_2_47_real = T1356 + T1354;
  assign T1354 = $signed(T1355) / $signed(22'h100000);
  assign T1355 = $signed(31'h29c4cf50) * $signed(16'h0);
  assign T1356 = $signed(T1357) / $signed(22'h100000);
  assign T1357 = $signed(31'h4f8253bf) * $signed(16'h1);
  assign T1358 = T383[1'h0:1'h0];
  assign T1359 = T383[1'h1:1'h1];
  assign T1360 = T383[2'h2:2'h2];
  assign T1361 = T383[2'h3:2'h3];
  assign T1362 = T1489 ? T1419 : T1363;
  assign T1363 = T1418 ? T1388 : T1364;
  assign T1364 = T1387 ? T1375 : T1365;
  assign T1365 = T1374 ? twiddle3_2_49_real : twiddle3_2_48_real;
  assign twiddle3_2_48_real = T1368 + T1366;
  assign T1366 = $signed(T1367) / $signed(22'h100000);
  assign T1367 = $signed(31'h2734d8ea) * $signed(16'h0);
  assign T1368 = $signed(T1369) / $signed(22'h100000);
  assign T1369 = $signed(31'h4d6a34de) * $signed(16'h1);
  assign twiddle3_2_49_real = T1372 + T1370;
  assign T1370 = $signed(T1371) / $signed(22'h100000);
  assign T1371 = $signed(31'h248a0caa) * $signed(16'h0);
  assign T1372 = $signed(T1373) / $signed(22'h100000);
  assign T1373 = $signed(31'h4b74b5a6) * $signed(16'h1);
  assign T1374 = T383[1'h0:1'h0];
  assign T1375 = T1386 ? twiddle3_2_51_real : twiddle3_2_50_real;
  assign twiddle3_2_50_real = T1378 + T1376;
  assign T1376 = $signed(T1377) / $signed(22'h100000);
  assign T1377 = $signed(31'h21c63de7) * $signed(16'h0);
  assign T1378 = $signed(T1379) / $signed(22'h100000);
  assign T1379 = $signed(31'h49a32d5a) * $signed(16'h1);
  assign twiddle3_2_51_real = T1384 + T1380;
  assign T1380 = {T1383, T1381};
  assign T1381 = $signed(T1382) / $signed(22'h100000);
  assign T1382 = $signed(30'h1eeb511b) * $signed(16'h0);
  assign T1383 = T1381[6'h2d:6'h2d];
  assign T1384 = $signed(T1385) / $signed(22'h100000);
  assign T1385 = $signed(31'h47f6da9c) * $signed(16'h1);
  assign T1386 = T383[1'h0:1'h0];
  assign T1387 = T383[1'h1:1'h1];
  assign T1388 = T1417 ? T1403 : T1389;
  assign T1389 = T1402 ? twiddle3_2_53_real : twiddle3_2_52_real;
  assign twiddle3_2_52_real = T1394 + T1390;
  assign T1390 = {T1393, T1391};
  assign T1391 = $signed(T1392) / $signed(22'h100000);
  assign T1392 = $signed(30'h1bfb3a90) * $signed(16'h0);
  assign T1393 = T1391[6'h2d:6'h2d];
  assign T1394 = $signed(T1395) / $signed(22'h100000);
  assign T1395 = $signed(31'h4670e29a) * $signed(16'h1);
  assign twiddle3_2_53_real = T1400 + T1396;
  assign T1396 = {T1399, T1397};
  assign T1397 = $signed(T1398) / $signed(22'h100000);
  assign T1398 = $signed(30'h18f7fd0d) * $signed(16'h0);
  assign T1399 = T1397[6'h2d:6'h2d];
  assign T1400 = $signed(T1401) / $signed(22'h100000);
  assign T1401 = $signed(31'h4512503e) * $signed(16'h1);
  assign T1402 = T383[1'h0:1'h0];
  assign T1403 = T1416 ? twiddle3_2_55_real : twiddle3_2_54_real;
  assign twiddle3_2_54_real = T1408 + T1404;
  assign T1404 = {T1407, T1405};
  assign T1405 = $signed(T1406) / $signed(22'h100000);
  assign T1406 = $signed(30'h15e3a874) * $signed(16'h0);
  assign T1407 = T1405[6'h2d:6'h2d];
  assign T1408 = $signed(T1409) / $signed(22'h100000);
  assign T1409 = $signed(31'h43dc137c) * $signed(16'h1);
  assign twiddle3_2_55_real = T1414 + T1410;
  assign T1410 = {T1413, T1411};
  assign T1411 = $signed(T1412) / $signed(22'h100000);
  assign T1412 = $signed(30'h12c0585b) * $signed(16'h0);
  assign T1413 = T1411[6'h2d:6'h2d];
  assign T1414 = $signed(T1415) / $signed(22'h100000);
  assign T1415 = $signed(31'h42cf00ad) * $signed(16'h1);
  assign T1416 = T383[1'h0:1'h0];
  assign T1417 = T383[1'h1:1'h1];
  assign T1418 = T383[2'h2:2'h2];
  assign T1419 = T1488 ? T1454 : T1420;
  assign T1420 = T1453 ? T1437 : T1421;
  assign T1421 = T1436 ? twiddle3_2_57_real : twiddle3_2_56_real;
  assign twiddle3_2_56_real = T1427 + T1422;
  assign T1422 = {T1425, T1423};
  assign T1423 = $signed(T1424) / $signed(22'h100000);
  assign T1424 = $signed(29'hf903299) * $signed(16'h0);
  assign T1425 = T1426 ? 2'h3 : 2'h0;
  assign T1426 = T1423[6'h2c:6'h2c];
  assign T1427 = $signed(T1428) / $signed(22'h100000);
  assign T1428 = $signed(31'h41ebcffd) * $signed(16'h1);
  assign twiddle3_2_57_real = T1434 + T1429;
  assign T1429 = {T1432, T1430};
  assign T1430 = $signed(T1431) / $signed(22'h100000);
  assign T1431 = $signed(29'hc5565ce) * $signed(16'h0);
  assign T1432 = T1433 ? 2'h3 : 2'h0;
  assign T1433 = T1430[6'h2c:6'h2c];
  assign T1434 = $signed(T1435) / $signed(22'h100000);
  assign T1435 = $signed(31'h41331ced) * $signed(16'h1);
  assign T1436 = T383[1'h0:1'h0];
  assign T1437 = T1452 ? twiddle3_2_59_real : twiddle3_2_58_real;
  assign twiddle3_2_58_real = T1443 + T1438;
  assign T1438 = {T1441, T1439};
  assign T1439 = $signed(T1440) / $signed(22'h100000);
  assign T1440 = $signed(29'h91227e2) * $signed(16'h0);
  assign T1441 = T1442 ? 2'h3 : 2'h0;
  assign T1442 = T1439[6'h2c:6'h2c];
  assign T1443 = $signed(T1444) / $signed(22'h100000);
  assign T1444 = $signed(31'h40a565e9) * $signed(16'h1);
  assign twiddle3_2_59_real = T1450 + T1445;
  assign T1445 = {T1448, T1446};
  assign T1446 = $signed(T1447) / $signed(22'h100000);
  assign T1447 = $signed(28'h5c8b488) * $signed(16'h0);
  assign T1448 = T1449 ? 3'h7 : 3'h0;
  assign T1449 = T1446[6'h2b:6'h2b];
  assign T1450 = $signed(T1451) / $signed(22'h100000);
  assign T1451 = $signed(31'h40430bef) * $signed(16'h1);
  assign T1452 = T383[1'h0:1'h0];
  assign T1453 = T383[1'h1:1'h1];
  assign T1454 = T1487 ? T1471 : T1455;
  assign T1455 = T1470 ? twiddle3_2_61_real : twiddle3_2_60_real;
  assign twiddle3_2_60_real = T1461 + T1456;
  assign T1456 = {T1459, T1457};
  assign T1457 = $signed(T1458) / $signed(22'h100000);
  assign T1458 = $signed(27'h27b4bb1) * $signed(16'h0);
  assign T1459 = T1460 ? 4'hf : 4'h0;
  assign T1460 = T1457[6'h2a:6'h2a];
  assign T1461 = $signed(T1462) / $signed(22'h100000);
  assign T1462 = $signed(31'h400c5251) * $signed(16'h1);
  assign twiddle3_2_61_real = T1468 + T1463;
  assign T1463 = {T1466, T1464};
  assign T1464 = $signed(T1465) / $signed(22'h100000);
  assign T1465 = $signed(25'h12c3005) * $signed(16'h0);
  assign T1466 = T1467 ? 6'h3f : 6'h0;
  assign T1467 = T1464[6'h28:6'h28];
  assign T1468 = $signed(T1469) / $signed(22'h100000);
  assign T1469 = $signed(31'h40015e85) * $signed(16'h1);
  assign T1470 = T383[1'h0:1'h0];
  assign T1471 = T1486 ? twiddle3_2_63_real : twiddle3_2_62_real;
  assign twiddle3_2_62_real = T1477 + T1472;
  assign T1472 = {T1475, T1473};
  assign T1473 = $signed(T1474) / $signed(22'h100000);
  assign T1474 = $signed(28'hbdda552) * $signed(16'h0);
  assign T1475 = T1476 ? 3'h7 : 3'h0;
  assign T1476 = T1473[6'h2b:6'h2b];
  assign T1477 = $signed(T1478) / $signed(22'h100000);
  assign T1478 = $signed(31'h4022380a) * $signed(16'h1);
  assign twiddle3_2_63_real = T1484 + T1479;
  assign T1479 = {T1482, T1480};
  assign T1480 = $signed(T1481) / $signed(22'h100000);
  assign T1481 = $signed(28'h891ef07) * $signed(16'h0);
  assign T1482 = T1483 ? 3'h7 : 3'h0;
  assign T1483 = T1480[6'h2b:6'h2b];
  assign T1484 = $signed(T1485) / $signed(22'h100000);
  assign T1485 = $signed(31'h406ec863) * $signed(16'h1);
  assign T1486 = T383[1'h0:1'h0];
  assign T1487 = T383[1'h1:1'h1];
  assign T1488 = T383[2'h2:2'h2];
  assign T1489 = T383[2'h3:2'h3];
  assign T1490 = T383[3'h4:3'h4];
  assign T1491 = T1245[6'h2e:6'h2e];
  assign T1492 = T383[3'h5:3'h5];
  assign T1493 = {T1610, T1494};
  assign T1494 = T1609 ? twiddle3_2_80_real : T1495;
  assign T1495 = T1604 ? T1558 : T1496;
  assign T1496 = T1557 ? T1529 : T1497;
  assign T1497 = T1528 ? T1514 : T1498;
  assign T1498 = T1513 ? twiddle3_2_65_real : twiddle3_2_64_real;
  assign twiddle3_2_64_real = T1504 + T1499;
  assign T1499 = {T1502, T1500};
  assign T1500 = $signed(T1501) / $signed(22'h100000);
  assign T1501 = $signed(29'h154b4ea1) * $signed(16'h0);
  assign T1502 = T1503 ? 2'h3 : 2'h0;
  assign T1503 = T1500[6'h2c:6'h2c];
  assign T1504 = $signed(T1505) / $signed(22'h100000);
  assign T1505 = $signed(31'h40e6db28) * $signed(16'h1);
  assign twiddle3_2_65_real = T1511 + T1506;
  assign T1506 = {T1509, T1507};
  assign T1507 = $signed(T1508) / $signed(22'h100000);
  assign T1508 = $signed(29'h120c0223) * $signed(16'h0);
  assign T1509 = T1510 ? 2'h3 : 2'h0;
  assign T1510 = T1507[6'h2c:6'h2c];
  assign T1511 = $signed(T1512) / $signed(22'h100000);
  assign T1512 = $signed(31'h418a1e2b) * $signed(16'h1);
  assign T1513 = T383[1'h0:1'h0];
  assign T1514 = T1527 ? twiddle3_2_67_real : twiddle3_2_66_real;
  assign twiddle3_2_66_real = T1519 + T1515;
  assign T1515 = {T1518, T1516};
  assign T1516 = $signed(T1517) / $signed(22'h100000);
  assign T1517 = $signed(30'h2ed6428a) * $signed(16'h0);
  assign T1518 = T1516[6'h2d:6'h2d];
  assign T1519 = $signed(T1520) / $signed(22'h100000);
  assign T1520 = $signed(31'h425821ac) * $signed(16'h1);
  assign twiddle3_2_67_real = T1525 + T1521;
  assign T1521 = {T1524, T1522};
  assign T1522 = $signed(T1523) / $signed(22'h100000);
  assign T1523 = $signed(30'h2bac424d) * $signed(16'h0);
  assign T1524 = T1522[6'h2d:6'h2d];
  assign T1525 = $signed(T1526) / $signed(22'h100000);
  assign T1526 = $signed(31'h435058a9) * $signed(16'h1);
  assign T1527 = T383[1'h0:1'h0];
  assign T1528 = T383[1'h1:1'h1];
  assign T1529 = T1556 ? T1544 : T1530;
  assign T1530 = T1543 ? twiddle3_2_69_real : twiddle3_2_68_real;
  assign twiddle3_2_68_real = T1535 + T1531;
  assign T1531 = {T1534, T1532};
  assign T1532 = $signed(T1533) / $signed(22'h100000);
  assign T1533 = $signed(30'h28902bd4) * $signed(16'h0);
  assign T1534 = T1532[6'h2d:6'h2d];
  assign T1535 = $signed(T1536) / $signed(22'h100000);
  assign T1536 = $signed(31'h4472193c) * $signed(16'h1);
  assign twiddle3_2_69_real = T1541 + T1537;
  assign T1537 = {T1540, T1538};
  assign T1538 = $signed(T1539) / $signed(22'h100000);
  assign T1539 = $signed(30'h25842006) * $signed(16'h0);
  assign T1540 = T1538[6'h2d:6'h2d];
  assign T1541 = $signed(T1542) / $signed(22'h100000);
  assign T1542 = $signed(31'h45bc9d14) * $signed(16'h1);
  assign T1543 = T383[1'h0:1'h0];
  assign T1544 = T1555 ? twiddle3_2_71_real : twiddle3_2_70_real;
  assign twiddle3_2_70_real = T1549 + T1545;
  assign T1545 = {T1548, T1546};
  assign T1546 = $signed(T1547) / $signed(22'h100000);
  assign T1547 = $signed(30'h228a34cc) * $signed(16'h0);
  assign T1548 = T1546[6'h2d:6'h2d];
  assign T1549 = $signed(T1550) / $signed(22'h100000);
  assign T1550 = $signed(31'h472f01f5) * $signed(16'h1);
  assign twiddle3_2_71_real = T1553 + T1551;
  assign T1551 = $signed(T1552) / $signed(22'h100000);
  assign T1552 = $signed(31'h5fa473a7) * $signed(16'h0);
  assign T1553 = $signed(T1554) / $signed(22'h100000);
  assign T1554 = $signed(31'h48c84a5b) * $signed(16'h1);
  assign T1555 = T383[1'h0:1'h0];
  assign T1556 = T383[1'h1:1'h1];
  assign T1557 = T383[2'h2:2'h2];
  assign T1558 = T1603 ? T1581 : T1559;
  assign T1559 = T1580 ? T1570 : T1560;
  assign T1560 = T1569 ? twiddle3_2_73_real : twiddle3_2_72_real;
  assign twiddle3_2_72_real = T1563 + T1561;
  assign T1561 = $signed(T1562) / $signed(22'h100000);
  assign T1562 = $signed(31'h5cd4d84c) * $signed(16'h0);
  assign T1563 = $signed(T1564) / $signed(22'h100000);
  assign T1564 = $signed(31'h4a875e22) * $signed(16'h1);
  assign twiddle3_2_73_real = T1567 + T1565;
  assign T1565 = $signed(T1566) / $signed(22'h100000);
  assign T1566 = $signed(31'h5a1d4f46) * $signed(16'h0);
  assign T1567 = $signed(T1568) / $signed(22'h100000);
  assign T1568 = $signed(31'h4c6b0b48) * $signed(16'h1);
  assign T1569 = T383[1'h0:1'h0];
  assign T1570 = T1579 ? twiddle3_2_75_real : twiddle3_2_74_real;
  assign twiddle3_2_74_real = T1573 + T1571;
  assign T1571 = $signed(T1572) / $signed(22'h100000);
  assign T1572 = $signed(31'h577fb4a6) * $signed(16'h0);
  assign T1573 = $signed(T1574) / $signed(22'h100000);
  assign T1574 = $signed(31'h4e7206bd) * $signed(16'h1);
  assign twiddle3_2_75_real = T1577 + T1575;
  assign T1575 = $signed(T1576) / $signed(22'h100000);
  assign T1576 = $signed(31'h54fdd2bf) * $signed(16'h0);
  assign T1577 = $signed(T1578) / $signed(22'h100000);
  assign T1578 = $signed(31'h509aed49) * $signed(16'h1);
  assign T1579 = T383[1'h0:1'h0];
  assign T1580 = T383[1'h1:1'h1];
  assign T1581 = T1602 ? T1592 : T1582;
  assign T1582 = T1591 ? twiddle3_2_77_real : twiddle3_2_76_real;
  assign twiddle3_2_76_real = T1585 + T1583;
  assign T1583 = $signed(T1584) / $signed(22'h100000);
  assign T1584 = $signed(31'h529960e8) * $signed(16'h0);
  assign T1585 = $signed(T1586) / $signed(22'h100000);
  assign T1586 = $signed(31'h52e4447b) * $signed(16'h1);
  assign twiddle3_2_77_real = T1589 + T1587;
  assign T1587 = $signed(T1588) / $signed(22'h100000);
  assign T1588 = $signed(31'h50540254) * $signed(16'h0);
  assign T1589 = $signed(T1590) / $signed(22'h100000);
  assign T1590 = $signed(31'h554c7bad) * $signed(16'h1);
  assign T1591 = T383[1'h0:1'h0];
  assign T1592 = T1601 ? twiddle3_2_79_real : twiddle3_2_78_real;
  assign twiddle3_2_78_real = T1595 + T1593;
  assign T1593 = $signed(T1594) / $signed(22'h100000);
  assign T1594 = $signed(31'h4e2f44f0) * $signed(16'h0);
  assign T1595 = $signed(T1596) / $signed(22'h100000);
  assign T1596 = $signed(31'h57d1ed19) * $signed(16'h1);
  assign twiddle3_2_79_real = T1599 + T1597;
  assign T1597 = $signed(T1598) / $signed(22'h100000);
  assign T1598 = $signed(31'h4c2ca054) * $signed(16'h0);
  assign T1599 = $signed(T1600) / $signed(22'h100000);
  assign T1600 = $signed(31'h5a72def6) * $signed(16'h1);
  assign T1601 = T383[1'h0:1'h0];
  assign T1602 = T383[1'h1:1'h1];
  assign T1603 = T383[2'h2:2'h2];
  assign T1604 = T383[2'h3:2'h3];
  assign twiddle3_2_80_real = T1607 + T1605;
  assign T1605 = $signed(T1606) / $signed(22'h100000);
  assign T1606 = $signed(31'h4a4d74c1) * $signed(16'h0);
  assign T1607 = $signed(T1608) / $signed(22'h100000);
  assign T1608 = $signed(31'h5d2d84aa) * $signed(16'h1);
  assign T1609 = T383[3'h4:3'h4];
  assign T1610 = T1494[6'h2e:6'h2e];
  assign T1611 = T383[3'h6:3'h6];
  assign io_t3_1out_imag = T1612;
  assign T1612 = T1613[4'hf:1'h0];
  assign T1613 = T2264 ? T2121 : T1614;
  assign T1614 = T2120 ? T1869 : T1615;
  assign T1615 = T1868 ? T1762 : T1616;
  assign T1616 = T1761 ? T1695 : T1617;
  assign T1617 = T1694 ? T1658 : T1618;
  assign T1618 = T1657 ? T1639 : T1619;
  assign T1619 = T1636 ? T1627 : twiddle3_1_0_imag;
  assign twiddle3_1_0_imag = T1625 + T1620;
  assign T1620 = {T1623, T1621};
  assign T1621 = $signed(T1622) / $signed(22'h100000);
  assign T1622 = $signed(1'h0) * $signed(16'hffff);
  assign T1623 = T1624 ? 31'h7fffffff : 31'h0;
  assign T1624 = T1621[5'h10:5'h10];
  assign T1625 = $signed(T1626) / $signed(22'h100000);
  assign T1626 = $signed(32'h40000000) * $signed(16'h0);
  assign T1627 = {T1635, twiddle3_1_1_imag};
  assign twiddle3_1_1_imag = T1633 + T1628;
  assign T1628 = {T1631, T1629};
  assign T1629 = $signed(T1630) / $signed(22'h100000);
  assign T1630 = $signed(26'h1a796e6) * $signed(16'hffff);
  assign T1631 = T1632 ? 5'h1f : 5'h0;
  assign T1632 = T1629[6'h29:6'h29];
  assign T1633 = $signed(T1634) / $signed(22'h100000);
  assign T1634 = $signed(31'h3ffa85fb) * $signed(16'h0);
  assign T1635 = twiddle3_1_1_imag[6'h2e:6'h2e];
  assign T1636 = T1637[1'h0:1'h0];
  assign T1637 = T1638;
  assign T1638 = io_in3[3'h6:1'h0];
  assign T1639 = {T1656, T1640};
  assign T1640 = T1655 ? twiddle3_1_3_imag : twiddle3_1_2_imag;
  assign twiddle3_1_2_imag = T1646 + T1641;
  assign T1641 = {T1644, T1642};
  assign T1642 = $signed(T1643) / $signed(22'h100000);
  assign T1643 = $signed(27'h34ee54e) * $signed(16'hffff);
  assign T1644 = T1645 ? 4'hf : 4'h0;
  assign T1645 = T1642[6'h2a:6'h2a];
  assign T1646 = $signed(T1647) / $signed(22'h100000);
  assign T1647 = $signed(31'h3fea18df) * $signed(16'h0);
  assign twiddle3_1_3_imag = T1653 + T1648;
  assign T1648 = {T1651, T1649};
  assign T1649 = $signed(T1650) / $signed(22'h100000);
  assign T1650 = $signed(28'h4f5a2c5) * $signed(16'hffff);
  assign T1651 = T1652 ? 3'h7 : 3'h0;
  assign T1652 = T1649[6'h2b:6'h2b];
  assign T1653 = $signed(T1654) / $signed(22'h100000);
  assign T1654 = $signed(31'h3fcebb7b) * $signed(16'h0);
  assign T1655 = T1637[1'h0:1'h0];
  assign T1656 = T1640[6'h2e:6'h2e];
  assign T1657 = T1637[1'h1:1'h1];
  assign T1658 = {T1693, T1659};
  assign T1659 = T1692 ? T1676 : T1660;
  assign T1660 = T1675 ? twiddle3_1_5_imag : twiddle3_1_4_imag;
  assign twiddle3_1_4_imag = T1666 + T1661;
  assign T1661 = {T1664, T1662};
  assign T1662 = $signed(T1663) / $signed(22'h100000);
  assign T1663 = $signed(28'h69b86f1) * $signed(16'hffff);
  assign T1664 = T1665 ? 3'h7 : 3'h0;
  assign T1665 = T1662[6'h2b:6'h2b];
  assign T1666 = $signed(T1667) / $signed(22'h100000);
  assign T1667 = $signed(31'h3fa8727d) * $signed(16'h0);
  assign twiddle3_1_5_imag = T1673 + T1668;
  assign T1668 = {T1671, T1669};
  assign T1669 = $signed(T1670) / $signed(22'h100000);
  assign T1670 = $signed(29'h840499e) * $signed(16'hffff);
  assign T1671 = T1672 ? 2'h3 : 2'h0;
  assign T1672 = T1669[6'h2c:6'h2c];
  assign T1673 = $signed(T1674) / $signed(22'h100000);
  assign T1674 = $signed(31'h3f774472) * $signed(16'h0);
  assign T1675 = T1637[1'h0:1'h0];
  assign T1676 = T1691 ? twiddle3_1_7_imag : twiddle3_1_6_imag;
  assign twiddle3_1_6_imag = T1682 + T1677;
  assign T1677 = {T1680, T1678};
  assign T1678 = $signed(T1679) / $signed(22'h100000);
  assign T1679 = $signed(29'h9e3a2ca) * $signed(16'hffff);
  assign T1680 = T1681 ? 2'h3 : 2'h0;
  assign T1681 = T1678[6'h2c:6'h2c];
  assign T1682 = $signed(T1683) / $signed(22'h100000);
  assign T1683 = $signed(31'h3f3b39c7) * $signed(16'h0);
  assign twiddle3_1_7_imag = T1689 + T1684;
  assign T1684 = {T1687, T1685};
  assign T1685 = $signed(T1686) / $signed(22'h100000);
  assign T1686 = $signed(29'hb854aaf) * $signed(16'hffff);
  assign T1687 = T1688 ? 2'h3 : 2'h0;
  assign T1688 = T1685[6'h2c:6'h2c];
  assign T1689 = $signed(T1690) / $signed(22'h100000);
  assign T1690 = $signed(31'h3ef45cc0) * $signed(16'h0);
  assign T1691 = T1637[1'h0:1'h0];
  assign T1692 = T1637[1'h1:1'h1];
  assign T1693 = T1659[6'h2e:6'h2e];
  assign T1694 = T1637[2'h2:2'h2];
  assign T1695 = {T1760, T1696};
  assign T1696 = T1759 ? T1729 : T1697;
  assign T1697 = T1728 ? T1714 : T1698;
  assign T1698 = T1713 ? twiddle3_1_9_imag : twiddle3_1_8_imag;
  assign twiddle3_1_8_imag = T1704 + T1699;
  assign T1699 = {T1702, T1700};
  assign T1700 = $signed(T1701) / $signed(22'h100000);
  assign T1701 = $signed(29'hd24f9d3) * $signed(16'hffff);
  assign T1702 = T1703 ? 2'h3 : 2'h0;
  assign T1703 = T1700[6'h2c:6'h2c];
  assign T1704 = $signed(T1705) / $signed(22'h100000);
  assign T1705 = $signed(31'h3ea2b980) * $signed(16'h0);
  assign twiddle3_1_9_imag = T1711 + T1706;
  assign T1706 = {T1709, T1707};
  assign T1707 = $signed(T1708) / $signed(22'h100000);
  assign T1708 = $signed(29'hec26911) * $signed(16'hffff);
  assign T1709 = T1710 ? 2'h3 : 2'h0;
  assign T1710 = T1707[6'h2c:6'h2c];
  assign T1711 = $signed(T1712) / $signed(22'h100000);
  assign T1712 = $signed(31'h3e465dfe) * $signed(16'h0);
  assign T1713 = T1637[1'h0:1'h0];
  assign T1714 = T1727 ? twiddle3_1_11_imag : twiddle3_1_10_imag;
  assign twiddle3_1_10_imag = T1719 + T1715;
  assign T1715 = {T1718, T1716};
  assign T1716 = $signed(T1717) / $signed(22'h100000);
  assign T1717 = $signed(30'h105d51a8) * $signed(16'hffff);
  assign T1718 = T1716[6'h2d:6'h2d];
  assign T1719 = $signed(T1720) / $signed(22'h100000);
  assign T1720 = $signed(31'h3ddf5a09) * $signed(16'h0);
  assign twiddle3_1_11_imag = T1725 + T1721;
  assign T1721 = {T1724, T1722};
  assign T1722 = $signed(T1723) / $signed(22'h100000);
  assign T1723 = $signed(30'h11f56d44) * $signed(16'hffff);
  assign T1724 = T1722[6'h2d:6'h2d];
  assign T1725 = $signed(T1726) / $signed(22'h100000);
  assign T1726 = $signed(31'h3d6dbf43) * $signed(16'h0);
  assign T1727 = T1637[1'h0:1'h0];
  assign T1728 = T1637[1'h1:1'h1];
  assign T1729 = T1758 ? T1744 : T1730;
  assign T1730 = T1743 ? twiddle3_1_13_imag : twiddle3_1_12_imag;
  assign twiddle3_1_12_imag = T1735 + T1731;
  assign T1731 = {T1734, T1732};
  assign T1732 = $signed(T1733) / $signed(22'h100000);
  assign T1733 = $signed(30'h138a760d) * $signed(16'hffff);
  assign T1734 = T1732[6'h2d:6'h2d];
  assign T1735 = $signed(T1736) / $signed(22'h100000);
  assign T1736 = $signed(31'h3cf1a11d) * $signed(16'h0);
  assign twiddle3_1_13_imag = T1741 + T1737;
  assign T1737 = {T1740, T1738};
  assign T1738 = $signed(T1739) / $signed(22'h100000);
  assign T1739 = $signed(30'h151c26b1) * $signed(16'hffff);
  assign T1740 = T1738[6'h2d:6'h2d];
  assign T1741 = $signed(T1742) / $signed(22'h100000);
  assign T1742 = $signed(31'h3c6b14d5) * $signed(16'h0);
  assign T1743 = T1637[1'h0:1'h0];
  assign T1744 = T1757 ? twiddle3_1_15_imag : twiddle3_1_14_imag;
  assign twiddle3_1_14_imag = T1749 + T1745;
  assign T1745 = {T1748, T1746};
  assign T1746 = $signed(T1747) / $signed(22'h100000);
  assign T1747 = $signed(30'h16aa3a72) * $signed(16'hffff);
  assign T1748 = T1746[6'h2d:6'h2d];
  assign T1749 = $signed(T1750) / $signed(22'h100000);
  assign T1750 = $signed(31'h3bda3171) * $signed(16'h0);
  assign twiddle3_1_15_imag = T1755 + T1751;
  assign T1751 = {T1754, T1752};
  assign T1752 = $signed(T1753) / $signed(22'h100000);
  assign T1753 = $signed(30'h18346d2d) * $signed(16'hffff);
  assign T1754 = T1752[6'h2d:6'h2d];
  assign T1755 = $signed(T1756) / $signed(22'h100000);
  assign T1756 = $signed(31'h3b3f0fbf) * $signed(16'h0);
  assign T1757 = T1637[1'h0:1'h0];
  assign T1758 = T1637[1'h1:1'h1];
  assign T1759 = T1637[2'h2:2'h2];
  assign T1760 = T1696[6'h2e:6'h2e];
  assign T1761 = T1637[2'h3:2'h3];
  assign T1762 = {T1867, T1763};
  assign T1763 = T1866 ? T1820 : T1764;
  assign T1764 = T1819 ? T1795 : T1765;
  assign T1765 = T1794 ? T1780 : T1766;
  assign T1766 = T1779 ? twiddle3_1_17_imag : twiddle3_1_16_imag;
  assign twiddle3_1_16_imag = T1771 + T1767;
  assign T1767 = {T1770, T1768};
  assign T1768 = $signed(T1769) / $signed(22'h100000);
  assign T1769 = $signed(30'h19ba7b6c) * $signed(16'hffff);
  assign T1770 = T1768[6'h2d:6'h2d];
  assign T1771 = $signed(T1772) / $signed(22'h100000);
  assign T1772 = $signed(31'h3a99ca4a) * $signed(16'h0);
  assign twiddle3_1_17_imag = T1777 + T1773;
  assign T1773 = {T1776, T1774};
  assign T1774 = $signed(T1775) / $signed(22'h100000);
  assign T1775 = $signed(30'h1b3c226e) * $signed(16'hffff);
  assign T1776 = T1774[6'h2d:6'h2d];
  assign T1777 = $signed(T1778) / $signed(22'h100000);
  assign T1778 = $signed(31'h39ea7d5c) * $signed(16'h0);
  assign T1779 = T1637[1'h0:1'h0];
  assign T1780 = T1793 ? twiddle3_1_19_imag : twiddle3_1_18_imag;
  assign twiddle3_1_18_imag = T1785 + T1781;
  assign T1781 = {T1784, T1782};
  assign T1782 = $signed(T1783) / $signed(22'h100000);
  assign T1783 = $signed(30'h1cb92032) * $signed(16'hffff);
  assign T1784 = T1782[6'h2d:6'h2d];
  assign T1785 = $signed(T1786) / $signed(22'h100000);
  assign T1786 = $signed(31'h393146f5) * $signed(16'h0);
  assign twiddle3_1_19_imag = T1791 + T1787;
  assign T1787 = {T1790, T1788};
  assign T1788 = $signed(T1789) / $signed(22'h100000);
  assign T1789 = $signed(30'h1e313383) * $signed(16'hffff);
  assign T1790 = T1788[6'h2d:6'h2d];
  assign T1791 = $signed(T1792) / $signed(22'h100000);
  assign T1792 = $signed(31'h386e46c7) * $signed(16'h0);
  assign T1793 = T1637[1'h0:1'h0];
  assign T1794 = T1637[1'h1:1'h1];
  assign T1795 = T1818 ? T1808 : T1796;
  assign T1796 = T1807 ? twiddle3_1_21_imag : twiddle3_1_20_imag;
  assign twiddle3_1_20_imag = T1801 + T1797;
  assign T1797 = {T1800, T1798};
  assign T1798 = $signed(T1799) / $signed(22'h100000);
  assign T1799 = $signed(30'h1fa41c05) * $signed(16'hffff);
  assign T1800 = T1798[6'h2d:6'h2d];
  assign T1801 = $signed(T1802) / $signed(22'h100000);
  assign T1802 = $signed(31'h37a19e34) * $signed(16'h0);
  assign twiddle3_1_21_imag = T1805 + T1803;
  assign T1803 = $signed(T1804) / $signed(22'h100000);
  assign T1804 = $signed(31'h21119a3d) * $signed(16'hffff);
  assign T1805 = $signed(T1806) / $signed(22'h100000);
  assign T1806 = $signed(31'h36cb7040) * $signed(16'h0);
  assign T1807 = T1637[1'h0:1'h0];
  assign T1808 = T1817 ? twiddle3_1_23_imag : twiddle3_1_22_imag;
  assign twiddle3_1_22_imag = T1811 + T1809;
  assign T1809 = $signed(T1810) / $signed(22'h100000);
  assign T1810 = $signed(31'h22796f9d) * $signed(16'hffff);
  assign T1811 = $signed(T1812) / $signed(22'h100000);
  assign T1812 = $signed(31'h35ebe194) * $signed(16'h0);
  assign twiddle3_1_23_imag = T1815 + T1813;
  assign T1813 = $signed(T1814) / $signed(22'h100000);
  assign T1814 = $signed(31'h23db5e91) * $signed(16'hffff);
  assign T1815 = $signed(T1816) / $signed(22'h100000);
  assign T1816 = $signed(31'h35031873) * $signed(16'h0);
  assign T1817 = T1637[1'h0:1'h0];
  assign T1818 = T1637[1'h1:1'h1];
  assign T1819 = T1637[2'h2:2'h2];
  assign T1820 = T1865 ? T1843 : T1821;
  assign T1821 = T1842 ? T1832 : T1822;
  assign T1822 = T1831 ? twiddle3_1_25_imag : twiddle3_1_24_imag;
  assign twiddle3_1_24_imag = T1825 + T1823;
  assign T1823 = $signed(T1824) / $signed(22'h100000);
  assign T1824 = $signed(31'h25372a85) * $signed(16'hffff);
  assign T1825 = $signed(T1826) / $signed(22'h100000);
  assign T1826 = $signed(31'h34113cb3) * $signed(16'h0);
  assign twiddle3_1_25_imag = T1829 + T1827;
  assign T1827 = $signed(T1828) / $signed(22'h100000);
  assign T1828 = $signed(31'h268c97f3) * $signed(16'hffff);
  assign T1829 = $signed(T1830) / $signed(22'h100000);
  assign T1830 = $signed(31'h331677ba) * $signed(16'h0);
  assign T1831 = T1637[1'h0:1'h0];
  assign T1832 = T1841 ? twiddle3_1_27_imag : twiddle3_1_26_imag;
  assign twiddle3_1_26_imag = T1835 + T1833;
  assign T1833 = $signed(T1834) / $signed(22'h100000);
  assign T1834 = $signed(31'h27db6c6d) * $signed(16'hffff);
  assign T1835 = $signed(T1836) / $signed(22'h100000);
  assign T1836 = $signed(31'h3212f472) * $signed(16'h0);
  assign twiddle3_1_27_imag = T1839 + T1837;
  assign T1837 = $signed(T1838) / $signed(22'h100000);
  assign T1838 = $signed(31'h29236ea4) * $signed(16'hffff);
  assign T1839 = $signed(T1840) / $signed(22'h100000);
  assign T1840 = $signed(31'h3106df45) * $signed(16'h0);
  assign T1841 = T1637[1'h0:1'h0];
  assign T1842 = T1637[1'h1:1'h1];
  assign T1843 = T1864 ? T1854 : T1844;
  assign T1844 = T1853 ? twiddle3_1_29_imag : twiddle3_1_28_imag;
  assign twiddle3_1_28_imag = T1847 + T1845;
  assign T1845 = $signed(T1846) / $signed(22'h100000);
  assign T1846 = $signed(31'h2a646676) * $signed(16'hffff);
  assign T1847 = $signed(T1848) / $signed(22'h100000);
  assign T1848 = $signed(31'h2ff26615) * $signed(16'h0);
  assign twiddle3_1_29_imag = T1851 + T1849;
  assign T1849 = $signed(T1850) / $signed(22'h100000);
  assign T1850 = $signed(31'h2b9e1cf3) * $signed(16'hffff);
  assign T1851 = $signed(T1852) / $signed(22'h100000);
  assign T1852 = $signed(31'h2ed5b833) * $signed(16'h0);
  assign T1853 = T1637[1'h0:1'h0];
  assign T1854 = T1863 ? twiddle3_1_31_imag : twiddle3_1_30_imag;
  assign twiddle3_1_30_imag = T1857 + T1855;
  assign T1855 = $signed(T1856) / $signed(22'h100000);
  assign T1856 = $signed(31'h2cd05c6c) * $signed(16'hffff);
  assign T1857 = $signed(T1858) / $signed(22'h100000);
  assign T1858 = $signed(31'h2db10657) * $signed(16'h0);
  assign twiddle3_1_31_imag = T1861 + T1859;
  assign T1859 = $signed(T1860) / $signed(22'h100000);
  assign T1860 = $signed(31'h2dfaf076) * $signed(16'hffff);
  assign T1861 = $signed(T1862) / $signed(22'h100000);
  assign T1862 = $signed(31'h2c848299) * $signed(16'h0);
  assign T1863 = T1637[1'h0:1'h0];
  assign T1864 = T1637[1'h1:1'h1];
  assign T1865 = T1637[2'h2:2'h2];
  assign T1866 = T1637[2'h3:2'h3];
  assign T1867 = T1763[6'h2e:6'h2e];
  assign T1868 = T1637[3'h4:3'h4];
  assign T1869 = {T2119, T1870};
  assign T1870 = T2118 ? T1979 : T1871;
  assign T1871 = T1978 ? T1918 : T1872;
  assign T1872 = T1917 ? T1895 : T1873;
  assign T1873 = T1894 ? T1884 : T1874;
  assign T1874 = T1883 ? twiddle3_1_33_imag : twiddle3_1_32_imag;
  assign twiddle3_1_32_imag = T1877 + T1875;
  assign T1875 = $signed(T1876) / $signed(22'h100000);
  assign T1876 = $signed(31'h2f1da5f8) * $signed(16'hffff);
  assign T1877 = $signed(T1878) / $signed(22'h100000);
  assign T1878 = $signed(31'h2b506069) * $signed(16'h0);
  assign twiddle3_1_33_imag = T1881 + T1879;
  assign T1879 = $signed(T1880) / $signed(22'h100000);
  assign T1880 = $signed(31'h30384b31) * $signed(16'hffff);
  assign T1881 = $signed(T1882) / $signed(22'h100000);
  assign T1882 = $signed(31'h2a14d481) * $signed(16'h0);
  assign T1883 = T1637[1'h0:1'h0];
  assign T1884 = T1893 ? twiddle3_1_35_imag : twiddle3_1_34_imag;
  assign twiddle3_1_34_imag = T1887 + T1885;
  assign T1885 = $signed(T1886) / $signed(22'h100000);
  assign T1886 = $signed(31'h314aafc2) * $signed(16'hffff);
  assign T1887 = $signed(T1888) / $signed(22'h100000);
  assign T1888 = $signed(31'h28d214e4) * $signed(16'h0);
  assign twiddle3_1_35_imag = T1891 + T1889;
  assign T1889 = $signed(T1890) / $signed(22'h100000);
  assign T1890 = $signed(31'h3254a4b4) * $signed(16'hffff);
  assign T1891 = $signed(T1892) / $signed(22'h100000);
  assign T1892 = $signed(31'h278858cd) * $signed(16'h0);
  assign T1893 = T1637[1'h0:1'h0];
  assign T1894 = T1637[1'h1:1'h1];
  assign T1895 = T1916 ? T1906 : T1896;
  assign T1896 = T1905 ? twiddle3_1_37_imag : twiddle3_1_36_imag;
  assign twiddle3_1_36_imag = T1899 + T1897;
  assign T1897 = $signed(T1898) / $signed(22'h100000);
  assign T1898 = $signed(31'h3355fc84) * $signed(16'hffff);
  assign T1899 = $signed(T1900) / $signed(22'h100000);
  assign T1900 = $signed(31'h2637d8ab) * $signed(16'h0);
  assign twiddle3_1_37_imag = T1903 + T1901;
  assign T1901 = $signed(T1902) / $signed(22'h100000);
  assign T1902 = $signed(31'h344e8b25) * $signed(16'hffff);
  assign T1903 = $signed(T1904) / $signed(22'h100000);
  assign T1904 = $signed(31'h24e0ce16) * $signed(16'h0);
  assign T1905 = T1637[1'h0:1'h0];
  assign T1906 = T1915 ? twiddle3_1_39_imag : twiddle3_1_38_imag;
  assign twiddle3_1_38_imag = T1909 + T1907;
  assign T1907 = $signed(T1908) / $signed(22'h100000);
  assign T1908 = $signed(31'h353e260f) * $signed(16'hffff);
  assign T1909 = $signed(T1910) / $signed(22'h100000);
  assign T1910 = $signed(31'h238373c3) * $signed(16'h0);
  assign twiddle3_1_39_imag = T1913 + T1911;
  assign T1911 = $signed(T1912) / $signed(22'h100000);
  assign T1912 = $signed(31'h3624a440) * $signed(16'hffff);
  assign T1913 = $signed(T1914) / $signed(22'h100000);
  assign T1914 = $signed(31'h2220057c) * $signed(16'h0);
  assign T1915 = T1637[1'h0:1'h0];
  assign T1916 = T1637[1'h1:1'h1];
  assign T1917 = T1637[2'h2:2'h2];
  assign T1918 = T1977 ? T1947 : T1919;
  assign T1919 = T1946 ? T1932 : T1920;
  assign T1920 = T1931 ? twiddle3_1_41_imag : twiddle3_1_40_imag;
  assign twiddle3_1_40_imag = T1923 + T1921;
  assign T1921 = $signed(T1922) / $signed(22'h100000);
  assign T1922 = $signed(31'h3701de44) * $signed(16'hffff);
  assign T1923 = $signed(T1924) / $signed(22'h100000);
  assign T1924 = $signed(31'h20b6c016) * $signed(16'h0);
  assign twiddle3_1_41_imag = T1927 + T1925;
  assign T1925 = $signed(T1926) / $signed(22'h100000);
  assign T1926 = $signed(31'h37d5ae3f) * $signed(16'hffff);
  assign T1927 = {T1930, T1928};
  assign T1928 = $signed(T1929) / $signed(22'h100000);
  assign T1929 = $signed(30'h1f47e165) * $signed(16'h0);
  assign T1930 = T1928[6'h2d:6'h2d];
  assign T1931 = T1637[1'h0:1'h0];
  assign T1932 = T1945 ? twiddle3_1_43_imag : twiddle3_1_42_imag;
  assign twiddle3_1_42_imag = T1935 + T1933;
  assign T1933 = $signed(T1934) / $signed(22'h100000);
  assign T1934 = $signed(31'h389feff1) * $signed(16'hffff);
  assign T1935 = {T1938, T1936};
  assign T1936 = $signed(T1937) / $signed(22'h100000);
  assign T1937 = $signed(30'h1dd3a832) * $signed(16'h0);
  assign T1938 = T1936[6'h2d:6'h2d];
  assign twiddle3_1_43_imag = T1941 + T1939;
  assign T1939 = $signed(T1940) / $signed(22'h100000);
  assign T1940 = $signed(31'h396080bd) * $signed(16'hffff);
  assign T1941 = {T1944, T1942};
  assign T1942 = $signed(T1943) / $signed(22'h100000);
  assign T1943 = $signed(30'h1c5a5433) * $signed(16'h0);
  assign T1944 = T1942[6'h2d:6'h2d];
  assign T1945 = T1637[1'h0:1'h0];
  assign T1946 = T1637[1'h1:1'h1];
  assign T1947 = T1976 ? T1962 : T1948;
  assign T1948 = T1961 ? twiddle3_1_45_imag : twiddle3_1_44_imag;
  assign twiddle3_1_44_imag = T1951 + T1949;
  assign T1949 = $signed(T1950) / $signed(22'h100000);
  assign T1950 = $signed(31'h3a173fae) * $signed(16'hffff);
  assign T1951 = {T1954, T1952};
  assign T1952 = $signed(T1953) / $signed(22'h100000);
  assign T1953 = $signed(30'h1adc25fb) * $signed(16'h0);
  assign T1954 = T1952[6'h2d:6'h2d];
  assign twiddle3_1_45_imag = T1957 + T1955;
  assign T1955 = $signed(T1956) / $signed(22'h100000);
  assign T1956 = $signed(31'h3ac40d7d) * $signed(16'hffff);
  assign T1957 = {T1960, T1958};
  assign T1958 = $signed(T1959) / $signed(22'h100000);
  assign T1959 = $signed(30'h19595ef2) * $signed(16'h0);
  assign T1960 = T1958[6'h2d:6'h2d];
  assign T1961 = T1637[1'h0:1'h0];
  assign T1962 = T1975 ? twiddle3_1_47_imag : twiddle3_1_46_imag;
  assign twiddle3_1_46_imag = T1965 + T1963;
  assign T1963 = $signed(T1964) / $signed(22'h100000);
  assign T1964 = $signed(31'h3b66cc97) * $signed(16'hffff);
  assign T1965 = {T1968, T1966};
  assign T1966 = $signed(T1967) / $signed(22'h100000);
  assign T1967 = $signed(30'h17d2414a) * $signed(16'h0);
  assign T1968 = T1966[6'h2d:6'h2d];
  assign twiddle3_1_47_imag = T1971 + T1969;
  assign T1969 = $signed(T1970) / $signed(22'h100000);
  assign T1970 = $signed(31'h3bff6121) * $signed(16'hffff);
  assign T1971 = {T1974, T1972};
  assign T1972 = $signed(T1973) / $signed(22'h100000);
  assign T1973 = $signed(30'h16470ff4) * $signed(16'h0);
  assign T1974 = T1972[6'h2d:6'h2d];
  assign T1975 = T1637[1'h0:1'h0];
  assign T1976 = T1637[1'h1:1'h1];
  assign T1977 = T1637[2'h2:2'h2];
  assign T1978 = T1637[2'h3:2'h3];
  assign T1979 = T2117 ? T2047 : T1980;
  assign T1980 = T2046 ? T2012 : T1981;
  assign T1981 = T2011 ? T1996 : T1982;
  assign T1982 = T1995 ? twiddle3_1_49_imag : twiddle3_1_48_imag;
  assign twiddle3_1_48_imag = T1985 + T1983;
  assign T1983 = $signed(T1984) / $signed(22'h100000);
  assign T1984 = $signed(31'h3c8db0ff) * $signed(16'hffff);
  assign T1985 = {T1988, T1986};
  assign T1986 = $signed(T1987) / $signed(22'h100000);
  assign T1987 = $signed(30'h14b80e91) * $signed(16'h0);
  assign T1988 = T1986[6'h2d:6'h2d];
  assign twiddle3_1_49_imag = T1991 + T1989;
  assign T1989 = $signed(T1990) / $signed(22'h100000);
  assign T1990 = $signed(31'h3d11a3d6) * $signed(16'hffff);
  assign T1991 = {T1994, T1992};
  assign T1992 = $signed(T1993) / $signed(22'h100000);
  assign T1993 = $signed(30'h1325816c) * $signed(16'h0);
  assign T1994 = T1992[6'h2d:6'h2d];
  assign T1995 = T1637[1'h0:1'h0];
  assign T1996 = T2010 ? twiddle3_1_51_imag : twiddle3_1_50_imag;
  assign twiddle3_1_50_imag = T1999 + T1997;
  assign T1997 = $signed(T1998) / $signed(22'h100000);
  assign T1998 = $signed(31'h3d8b2310) * $signed(16'hffff);
  assign T1999 = {T2002, T2000};
  assign T2000 = $signed(T2001) / $signed(22'h100000);
  assign T2001 = $signed(30'h118fad69) * $signed(16'h0);
  assign T2002 = T2000[6'h2d:6'h2d];
  assign twiddle3_1_51_imag = T2005 + T2003;
  assign T2003 = $signed(T2004) / $signed(22'h100000);
  assign T2004 = $signed(31'h3dfa19e2) * $signed(16'hffff);
  assign T2005 = {T2008, T2006};
  assign T2006 = $signed(T2007) / $signed(22'h100000);
  assign T2007 = $signed(29'hff6d7fd) * $signed(16'h0);
  assign T2008 = T2009 ? 2'h3 : 2'h0;
  assign T2009 = T2006[6'h2c:6'h2c];
  assign T2010 = T1637[1'h0:1'h0];
  assign T2011 = T1637[1'h1:1'h1];
  assign T2012 = T2045 ? T2029 : T2013;
  assign T2013 = T2028 ? twiddle3_1_53_imag : twiddle3_1_52_imag;
  assign twiddle3_1_52_imag = T2016 + T2014;
  assign T2014 = $signed(T2015) / $signed(22'h100000);
  assign T2015 = $signed(31'h3e5e754f) * $signed(16'hffff);
  assign T2016 = {T2019, T2017};
  assign T2017 = $signed(T2018) / $signed(22'h100000);
  assign T2018 = $signed(29'he5b4720) * $signed(16'h0);
  assign T2019 = T2020 ? 2'h3 : 2'h0;
  assign T2020 = T2017[6'h2c:6'h2c];
  assign twiddle3_1_53_imag = T2023 + T2021;
  assign T2021 = $signed(T2022) / $signed(22'h100000);
  assign T2022 = $signed(31'h3eb8242a) * $signed(16'hffff);
  assign T2023 = {T2026, T2024};
  assign T2024 = $signed(T2025) / $signed(22'h100000);
  assign T2025 = $signed(29'hcbd4142) * $signed(16'h0);
  assign T2026 = T2027 ? 2'h3 : 2'h0;
  assign T2027 = T2024[6'h2c:6'h2c];
  assign T2028 = T1637[1'h0:1'h0];
  assign T2029 = T2044 ? twiddle3_1_55_imag : twiddle3_1_54_imag;
  assign twiddle3_1_54_imag = T2032 + T2030;
  assign T2030 = $signed(T2031) / $signed(22'h100000);
  assign T2031 = $signed(31'h3f071719) * $signed(16'hffff);
  assign T2032 = {T2035, T2033};
  assign T2033 = $signed(T2034) / $signed(22'h100000);
  assign T2034 = $signed(29'hb1d0d3f) * $signed(16'h0);
  assign T2035 = T2036 ? 2'h3 : 2'h0;
  assign T2036 = T2033[6'h2c:6'h2c];
  assign twiddle3_1_55_imag = T2039 + T2037;
  assign T2037 = $signed(T2038) / $signed(22'h100000);
  assign T2038 = $signed(31'h3f4b4099) * $signed(16'hffff);
  assign T2039 = {T2042, T2040};
  assign T2040 = $signed(T2041) / $signed(22'h100000);
  assign T2041 = $signed(29'h97af251) * $signed(16'h0);
  assign T2042 = T2043 ? 2'h3 : 2'h0;
  assign T2043 = T2040[6'h2c:6'h2c];
  assign T2044 = T1637[1'h0:1'h0];
  assign T2045 = T1637[1'h1:1'h1];
  assign T2046 = T1637[2'h2:2'h2];
  assign T2047 = T2116 ? T2082 : T2048;
  assign T2048 = T2081 ? T2065 : T2049;
  assign T2049 = T2064 ? twiddle3_1_57_imag : twiddle3_1_56_imag;
  assign twiddle3_1_56_imag = T2052 + T2050;
  assign T2050 = $signed(T2051) / $signed(22'h100000);
  assign T2051 = $signed(31'h3f849500) * $signed(16'hffff);
  assign T2052 = {T2055, T2053};
  assign T2053 = $signed(T2054) / $signed(22'h100000);
  assign T2054 = $signed(28'h7d73808) * $signed(16'h0);
  assign T2055 = T2056 ? 3'h7 : 3'h0;
  assign T2056 = T2053[6'h2b:6'h2b];
  assign twiddle3_1_57_imag = T2059 + T2057;
  assign T2057 = $signed(T2058) / $signed(22'h100000);
  assign T2058 = $signed(31'h3fb30a7f) * $signed(16'hffff);
  assign T2059 = {T2062, T2060};
  assign T2060 = $signed(T2061) / $signed(22'h100000);
  assign T2061 = $signed(28'h6322638) * $signed(16'h0);
  assign T2062 = T2063 ? 3'h7 : 3'h0;
  assign T2063 = T2060[6'h2b:6'h2b];
  assign T2064 = T1637[1'h0:1'h0];
  assign T2065 = T2080 ? twiddle3_1_59_imag : twiddle3_1_58_imag;
  assign twiddle3_1_58_imag = T2068 + T2066;
  assign T2066 = $signed(T2067) / $signed(22'h100000);
  assign T2067 = $signed(31'h3fd69921) * $signed(16'hffff);
  assign T2068 = {T2071, T2069};
  assign T2069 = $signed(T2070) / $signed(22'h100000);
  assign T2070 = $signed(28'h48c04f3) * $signed(16'h0);
  assign T2071 = T2072 ? 3'h7 : 3'h0;
  assign T2072 = T2069[6'h2b:6'h2b];
  assign twiddle3_1_59_imag = T2075 + T2073;
  assign T2073 = $signed(T2074) / $signed(22'h100000);
  assign T2074 = $signed(31'h3fef3ad1) * $signed(16'hffff);
  assign T2075 = {T2078, T2076};
  assign T2076 = $signed(T2077) / $signed(22'h100000);
  assign T2077 = $signed(27'h2e51c76) * $signed(16'h0);
  assign T2078 = T2079 ? 4'hf : 4'h0;
  assign T2079 = T2076[6'h2a:6'h2a];
  assign T2080 = T1637[1'h0:1'h0];
  assign T2081 = T1637[1'h1:1'h1];
  assign T2082 = T2115 ? T2099 : T2083;
  assign T2083 = T2098 ? twiddle3_1_61_imag : twiddle3_1_60_imag;
  assign twiddle3_1_60_imag = T2086 + T2084;
  assign T2084 = $signed(T2085) / $signed(22'h100000);
  assign T2085 = $signed(31'h3ffceb58) * $signed(16'hffff);
  assign T2086 = {T2089, T2087};
  assign T2087 = $signed(T2088) / $signed(22'h100000);
  assign T2088 = $signed(26'h13db523) * $signed(16'h0);
  assign T2089 = T2090 ? 5'h1f : 5'h0;
  assign T2090 = T2087[6'h29:6'h29];
  assign twiddle3_1_61_imag = T2093 + T2091;
  assign T2091 = $signed(T2092) / $signed(22'h100000);
  assign T2092 = $signed(31'h3fffa85e) * $signed(16'hffff);
  assign T2093 = {T2096, T2094};
  assign T2094 = $signed(T2095) / $signed(22'h100000);
  assign T2095 = $signed(24'h961772) * $signed(16'h0);
  assign T2096 = T2097 ? 7'h7f : 7'h0;
  assign T2097 = T2094[6'h27:6'h27];
  assign T2098 = T1637[1'h0:1'h0];
  assign T2099 = T2114 ? twiddle3_1_63_imag : twiddle3_1_62_imag;
  assign twiddle3_1_62_imag = T2102 + T2100;
  assign T2100 = $signed(T2101) / $signed(22'h100000);
  assign T2101 = $signed(31'h3ff7716b) * $signed(16'hffff);
  assign T2102 = {T2105, T2103};
  assign T2103 = $signed(T2104) / $signed(22'h100000);
  assign T2104 = $signed(27'h5ee8bdf) * $signed(16'h0);
  assign T2105 = T2106 ? 4'hf : 4'h0;
  assign T2106 = T2103[6'h2a:6'h2a];
  assign twiddle3_1_63_imag = T2109 + T2107;
  assign T2107 = $signed(T2108) / $signed(22'h100000);
  assign T2108 = $signed(31'h3fe447e6) * $signed(16'hffff);
  assign T2109 = {T2112, T2110};
  assign T2110 = $signed(T2111) / $signed(22'h100000);
  assign T2111 = $signed(27'h4475aea) * $signed(16'h0);
  assign T2112 = T2113 ? 4'hf : 4'h0;
  assign T2113 = T2110[6'h2a:6'h2a];
  assign T2114 = T1637[1'h0:1'h0];
  assign T2115 = T1637[1'h1:1'h1];
  assign T2116 = T1637[2'h2:2'h2];
  assign T2117 = T1637[2'h3:2'h3];
  assign T2118 = T1637[3'h4:3'h4];
  assign T2119 = T1870[6'h2e:6'h2e];
  assign T2120 = T1637[3'h5:3'h5];
  assign T2121 = {T2263, T2122};
  assign T2122 = T2262 ? twiddle3_1_80_imag : T2123;
  assign T2123 = T2255 ? T2193 : T2124;
  assign T2124 = T2192 ? T2159 : T2125;
  assign T2125 = T2158 ? T2142 : T2126;
  assign T2126 = T2141 ? twiddle3_1_65_imag : twiddle3_1_64_imag;
  assign twiddle3_1_64_imag = T2129 + T2127;
  assign T2127 = $signed(T2128) / $signed(22'h100000);
  assign T2128 = $signed(31'h3fc62f18) * $signed(16'hffff);
  assign T2129 = {T2132, T2130};
  assign T2130 = $signed(T2131) / $signed(22'h100000);
  assign T2131 = $signed(28'haa0ccff) * $signed(16'h0);
  assign T2132 = T2133 ? 3'h7 : 3'h0;
  assign T2133 = T2130[6'h2b:6'h2b];
  assign twiddle3_1_65_imag = T2136 + T2134;
  assign T2134 = $signed(T2135) / $signed(22'h100000);
  assign T2135 = $signed(31'h3f9d2c27) * $signed(16'hffff);
  assign T2136 = {T2139, T2137};
  assign T2137 = $signed(T2138) / $signed(22'h100000);
  assign T2138 = $signed(28'h8fb2a6f) * $signed(16'h0);
  assign T2139 = T2140 ? 3'h7 : 3'h0;
  assign T2140 = T2137[6'h2b:6'h2b];
  assign T2141 = T1637[1'h0:1'h0];
  assign T2142 = T2157 ? twiddle3_1_67_imag : twiddle3_1_66_imag;
  assign twiddle3_1_66_imag = T2145 + T2143;
  assign T2143 = $signed(T2144) / $signed(22'h100000);
  assign T2144 = $signed(31'h3f694618) * $signed(16'hffff);
  assign T2145 = {T2148, T2146};
  assign T2146 = $signed(T2147) / $signed(22'h100000);
  assign T2147 = $signed(29'h1756bb64) * $signed(16'h0);
  assign T2148 = T2149 ? 2'h3 : 2'h0;
  assign T2149 = T2146[6'h2c:6'h2c];
  assign twiddle3_1_67_imag = T2152 + T2150;
  assign T2150 = $signed(T2151) / $signed(22'h100000);
  assign T2151 = $signed(31'h3f2a85cc) * $signed(16'hffff);
  assign T2152 = {T2155, T2153};
  assign T2153 = $signed(T2154) / $signed(22'h100000);
  assign T2154 = $signed(29'h15b3c7d2) * $signed(16'h0);
  assign T2155 = T2156 ? 2'h3 : 2'h0;
  assign T2156 = T2153[6'h2c:6'h2c];
  assign T2157 = T1637[1'h0:1'h0];
  assign T2158 = T1637[1'h1:1'h1];
  assign T2159 = T2191 ? T2176 : T2160;
  assign T2160 = T2175 ? twiddle3_1_69_imag : twiddle3_1_68_imag;
  assign twiddle3_1_68_imag = T2163 + T2161;
  assign T2161 = $signed(T2162) / $signed(22'h100000);
  assign T2162 = $signed(31'h3ee0f602) * $signed(16'hffff);
  assign T2163 = {T2166, T2164};
  assign T2164 = $signed(T2165) / $signed(22'h100000);
  assign T2165 = $signed(29'h1412976d) * $signed(16'h0);
  assign T2166 = T2167 ? 2'h3 : 2'h0;
  assign T2167 = T2164[6'h2c:6'h2c];
  assign twiddle3_1_69_imag = T2170 + T2168;
  assign T2168 = $signed(T2169) / $signed(22'h100000);
  assign T2169 = $signed(31'h3e8ca34f) * $signed(16'hffff);
  assign T2170 = {T2173, T2171};
  assign T2171 = $signed(T2172) / $signed(22'h100000);
  assign T2172 = $signed(29'h1273719b) * $signed(16'h0);
  assign T2173 = T2174 ? 2'h3 : 2'h0;
  assign T2174 = T2171[6'h2c:6'h2c];
  assign T2175 = T1637[1'h0:1'h0];
  assign T2176 = T2190 ? twiddle3_1_71_imag : twiddle3_1_70_imag;
  assign twiddle3_1_70_imag = T2179 + T2177;
  assign T2177 = $signed(T2178) / $signed(22'h100000);
  assign T2178 = $signed(31'h3e2d9c23) * $signed(16'hffff);
  assign T2179 = {T2182, T2180};
  assign T2180 = $signed(T2181) / $signed(22'h100000);
  assign T2181 = $signed(29'h10d69d68) * $signed(16'h0);
  assign T2182 = T2183 ? 2'h3 : 2'h0;
  assign T2183 = T2180[6'h2c:6'h2c];
  assign twiddle3_1_71_imag = T2186 + T2184;
  assign T2184 = $signed(T2185) / $signed(22'h100000);
  assign T2185 = $signed(31'h3dc3f0c1) * $signed(16'hffff);
  assign T2186 = {T2189, T2187};
  assign T2187 = $signed(T2188) / $signed(22'h100000);
  assign T2188 = $signed(30'h2f3c617d) * $signed(16'h0);
  assign T2189 = T2187[6'h2d:6'h2d];
  assign T2190 = T1637[1'h0:1'h0];
  assign T2191 = T1637[1'h1:1'h1];
  assign T2192 = T1637[2'h2:2'h2];
  assign T2193 = T2254 ? T2224 : T2194;
  assign T2194 = T2223 ? T2209 : T2195;
  assign T2195 = T2208 ? twiddle3_1_73_imag : twiddle3_1_72_imag;
  assign twiddle3_1_72_imag = T2198 + T2196;
  assign T2196 = $signed(T2197) / $signed(22'h100000);
  assign T2197 = $signed(31'h3d4fb33e) * $signed(16'hffff);
  assign T2198 = {T2201, T2199};
  assign T2199 = $signed(T2200) / $signed(22'h100000);
  assign T2200 = $signed(30'h2da5040e) * $signed(16'h0);
  assign T2201 = T2199[6'h2d:6'h2d];
  assign twiddle3_1_73_imag = T2204 + T2202;
  assign T2202 = $signed(T2203) / $signed(22'h100000);
  assign T2203 = $signed(31'h3cd0f77f) * $signed(16'hffff);
  assign T2204 = {T2207, T2205};
  assign T2205 = $signed(T2206) / $signed(22'h100000);
  assign T2206 = $signed(30'h2c10cad4) * $signed(16'h0);
  assign T2207 = T2205[6'h2d:6'h2d];
  assign T2208 = T1637[1'h0:1'h0];
  assign T2209 = T2222 ? twiddle3_1_75_imag : twiddle3_1_74_imag;
  assign twiddle3_1_74_imag = T2212 + T2210;
  assign T2210 = $signed(T2211) / $signed(22'h100000);
  assign T2211 = $signed(31'h3c47d336) * $signed(16'hffff);
  assign T2212 = {T2215, T2213};
  assign T2213 = $signed(T2214) / $signed(22'h100000);
  assign T2214 = $signed(30'h2a7ffafd) * $signed(16'h0);
  assign T2215 = T2213[6'h2d:6'h2d];
  assign twiddle3_1_75_imag = T2218 + T2216;
  assign T2216 = $signed(T2217) / $signed(22'h100000);
  assign T2217 = $signed(31'h3bb45dda) * $signed(16'hffff);
  assign T2218 = {T2221, T2219};
  assign T2219 = $signed(T2220) / $signed(22'h100000);
  assign T2220 = $signed(30'h28f2d921) * $signed(16'h0);
  assign T2221 = T2219[6'h2d:6'h2d];
  assign T2222 = T1637[1'h0:1'h0];
  assign T2223 = T1637[1'h1:1'h1];
  assign T2224 = T2253 ? T2239 : T2225;
  assign T2225 = T2238 ? twiddle3_1_77_imag : twiddle3_1_76_imag;
  assign twiddle3_1_76_imag = T2228 + T2226;
  assign T2226 = $signed(T2227) / $signed(22'h100000);
  assign T2227 = $signed(31'h3b16b0a8) * $signed(16'hffff);
  assign T2228 = {T2231, T2229};
  assign T2229 = $signed(T2230) / $signed(22'h100000);
  assign T2230 = $signed(30'h2769a939) * $signed(16'h0);
  assign T2231 = T2229[6'h2d:6'h2d];
  assign twiddle3_1_77_imag = T2234 + T2232;
  assign T2232 = $signed(T2233) / $signed(22'h100000);
  assign T2233 = $signed(31'h3a6ee69d) * $signed(16'hffff);
  assign T2234 = {T2237, T2235};
  assign T2235 = $signed(T2236) / $signed(22'h100000);
  assign T2236 = $signed(30'h25e4ae8e) * $signed(16'h0);
  assign T2237 = T2235[6'h2d:6'h2d];
  assign T2238 = T1637[1'h0:1'h0];
  assign T2239 = T2252 ? twiddle3_1_79_imag : twiddle3_1_78_imag;
  assign twiddle3_1_78_imag = T2242 + T2240;
  assign T2240 = $signed(T2241) / $signed(22'h100000);
  assign T2241 = $signed(31'h39bd1c70) * $signed(16'hffff);
  assign T2242 = {T2245, T2243};
  assign T2243 = $signed(T2244) / $signed(22'h100000);
  assign T2244 = $signed(30'h24642bb3) * $signed(16'h0);
  assign T2245 = T2243[6'h2d:6'h2d];
  assign twiddle3_1_79_imag = T2248 + T2246;
  assign T2246 = $signed(T2247) / $signed(22'h100000);
  assign T2247 = $signed(31'h3901708e) * $signed(16'hffff);
  assign T2248 = {T2251, T2249};
  assign T2249 = $signed(T2250) / $signed(22'h100000);
  assign T2250 = $signed(30'h22e86278) * $signed(16'h0);
  assign T2251 = T2249[6'h2d:6'h2d];
  assign T2252 = T1637[1'h0:1'h0];
  assign T2253 = T1637[1'h1:1'h1];
  assign T2254 = T1637[2'h2:2'h2];
  assign T2255 = T1637[2'h3:2'h3];
  assign twiddle3_1_80_imag = T2258 + T2256;
  assign T2256 = $signed(T2257) / $signed(22'h100000);
  assign T2257 = $signed(31'h383c0315) * $signed(16'hffff);
  assign T2258 = {T2261, T2259};
  assign T2259 = $signed(T2260) / $signed(22'h100000);
  assign T2260 = $signed(30'h217193da) * $signed(16'h0);
  assign T2261 = T2259[6'h2d:6'h2d];
  assign T2262 = T1637[3'h4:3'h4];
  assign T2263 = T2122[6'h2e:6'h2e];
  assign T2264 = T1637[3'h6:3'h6];
  assign io_t3_1out_real = T2265;
  assign T2265 = T2266[4'hf:1'h0];
  assign T2266 = T2915 ? T2772 : T2267;
  assign T2267 = T2771 ? T2520 : T2268;
  assign T2268 = T2519 ? T2413 : T2269;
  assign T2269 = T2412 ? T2346 : T2270;
  assign T2270 = T2345 ? T2309 : T2271;
  assign T2271 = T2308 ? T2290 : T2272;
  assign T2272 = T2289 ? T2280 : twiddle3_1_0_real;
  assign twiddle3_1_0_real = T2278 + T2273;
  assign T2273 = {T2276, T2274};
  assign T2274 = $signed(T2275) / $signed(22'h100000);
  assign T2275 = $signed(1'h0) * $signed(16'h0);
  assign T2276 = T2277 ? 31'h7fffffff : 31'h0;
  assign T2277 = T2274[5'h10:5'h10];
  assign T2278 = $signed(T2279) / $signed(22'h100000);
  assign T2279 = $signed(32'h40000000) * $signed(16'h1);
  assign T2280 = {T2288, twiddle3_1_1_real};
  assign twiddle3_1_1_real = T2286 + T2281;
  assign T2281 = {T2284, T2282};
  assign T2282 = $signed(T2283) / $signed(22'h100000);
  assign T2283 = $signed(26'h1a796e6) * $signed(16'h0);
  assign T2284 = T2285 ? 5'h1f : 5'h0;
  assign T2285 = T2282[6'h29:6'h29];
  assign T2286 = $signed(T2287) / $signed(22'h100000);
  assign T2287 = $signed(31'h3ffa85fb) * $signed(16'h1);
  assign T2288 = twiddle3_1_1_real[6'h2e:6'h2e];
  assign T2289 = T1637[1'h0:1'h0];
  assign T2290 = {T2307, T2291};
  assign T2291 = T2306 ? twiddle3_1_3_real : twiddle3_1_2_real;
  assign twiddle3_1_2_real = T2297 + T2292;
  assign T2292 = {T2295, T2293};
  assign T2293 = $signed(T2294) / $signed(22'h100000);
  assign T2294 = $signed(27'h34ee54e) * $signed(16'h0);
  assign T2295 = T2296 ? 4'hf : 4'h0;
  assign T2296 = T2293[6'h2a:6'h2a];
  assign T2297 = $signed(T2298) / $signed(22'h100000);
  assign T2298 = $signed(31'h3fea18df) * $signed(16'h1);
  assign twiddle3_1_3_real = T2304 + T2299;
  assign T2299 = {T2302, T2300};
  assign T2300 = $signed(T2301) / $signed(22'h100000);
  assign T2301 = $signed(28'h4f5a2c5) * $signed(16'h0);
  assign T2302 = T2303 ? 3'h7 : 3'h0;
  assign T2303 = T2300[6'h2b:6'h2b];
  assign T2304 = $signed(T2305) / $signed(22'h100000);
  assign T2305 = $signed(31'h3fcebb7b) * $signed(16'h1);
  assign T2306 = T1637[1'h0:1'h0];
  assign T2307 = T2291[6'h2e:6'h2e];
  assign T2308 = T1637[1'h1:1'h1];
  assign T2309 = {T2344, T2310};
  assign T2310 = T2343 ? T2327 : T2311;
  assign T2311 = T2326 ? twiddle3_1_5_real : twiddle3_1_4_real;
  assign twiddle3_1_4_real = T2317 + T2312;
  assign T2312 = {T2315, T2313};
  assign T2313 = $signed(T2314) / $signed(22'h100000);
  assign T2314 = $signed(28'h69b86f1) * $signed(16'h0);
  assign T2315 = T2316 ? 3'h7 : 3'h0;
  assign T2316 = T2313[6'h2b:6'h2b];
  assign T2317 = $signed(T2318) / $signed(22'h100000);
  assign T2318 = $signed(31'h3fa8727d) * $signed(16'h1);
  assign twiddle3_1_5_real = T2324 + T2319;
  assign T2319 = {T2322, T2320};
  assign T2320 = $signed(T2321) / $signed(22'h100000);
  assign T2321 = $signed(29'h840499e) * $signed(16'h0);
  assign T2322 = T2323 ? 2'h3 : 2'h0;
  assign T2323 = T2320[6'h2c:6'h2c];
  assign T2324 = $signed(T2325) / $signed(22'h100000);
  assign T2325 = $signed(31'h3f774472) * $signed(16'h1);
  assign T2326 = T1637[1'h0:1'h0];
  assign T2327 = T2342 ? twiddle3_1_7_real : twiddle3_1_6_real;
  assign twiddle3_1_6_real = T2333 + T2328;
  assign T2328 = {T2331, T2329};
  assign T2329 = $signed(T2330) / $signed(22'h100000);
  assign T2330 = $signed(29'h9e3a2ca) * $signed(16'h0);
  assign T2331 = T2332 ? 2'h3 : 2'h0;
  assign T2332 = T2329[6'h2c:6'h2c];
  assign T2333 = $signed(T2334) / $signed(22'h100000);
  assign T2334 = $signed(31'h3f3b39c7) * $signed(16'h1);
  assign twiddle3_1_7_real = T2340 + T2335;
  assign T2335 = {T2338, T2336};
  assign T2336 = $signed(T2337) / $signed(22'h100000);
  assign T2337 = $signed(29'hb854aaf) * $signed(16'h0);
  assign T2338 = T2339 ? 2'h3 : 2'h0;
  assign T2339 = T2336[6'h2c:6'h2c];
  assign T2340 = $signed(T2341) / $signed(22'h100000);
  assign T2341 = $signed(31'h3ef45cc0) * $signed(16'h1);
  assign T2342 = T1637[1'h0:1'h0];
  assign T2343 = T1637[1'h1:1'h1];
  assign T2344 = T2310[6'h2e:6'h2e];
  assign T2345 = T1637[2'h2:2'h2];
  assign T2346 = {T2411, T2347};
  assign T2347 = T2410 ? T2380 : T2348;
  assign T2348 = T2379 ? T2365 : T2349;
  assign T2349 = T2364 ? twiddle3_1_9_real : twiddle3_1_8_real;
  assign twiddle3_1_8_real = T2355 + T2350;
  assign T2350 = {T2353, T2351};
  assign T2351 = $signed(T2352) / $signed(22'h100000);
  assign T2352 = $signed(29'hd24f9d3) * $signed(16'h0);
  assign T2353 = T2354 ? 2'h3 : 2'h0;
  assign T2354 = T2351[6'h2c:6'h2c];
  assign T2355 = $signed(T2356) / $signed(22'h100000);
  assign T2356 = $signed(31'h3ea2b980) * $signed(16'h1);
  assign twiddle3_1_9_real = T2362 + T2357;
  assign T2357 = {T2360, T2358};
  assign T2358 = $signed(T2359) / $signed(22'h100000);
  assign T2359 = $signed(29'hec26911) * $signed(16'h0);
  assign T2360 = T2361 ? 2'h3 : 2'h0;
  assign T2361 = T2358[6'h2c:6'h2c];
  assign T2362 = $signed(T2363) / $signed(22'h100000);
  assign T2363 = $signed(31'h3e465dfe) * $signed(16'h1);
  assign T2364 = T1637[1'h0:1'h0];
  assign T2365 = T2378 ? twiddle3_1_11_real : twiddle3_1_10_real;
  assign twiddle3_1_10_real = T2370 + T2366;
  assign T2366 = {T2369, T2367};
  assign T2367 = $signed(T2368) / $signed(22'h100000);
  assign T2368 = $signed(30'h105d51a8) * $signed(16'h0);
  assign T2369 = T2367[6'h2d:6'h2d];
  assign T2370 = $signed(T2371) / $signed(22'h100000);
  assign T2371 = $signed(31'h3ddf5a09) * $signed(16'h1);
  assign twiddle3_1_11_real = T2376 + T2372;
  assign T2372 = {T2375, T2373};
  assign T2373 = $signed(T2374) / $signed(22'h100000);
  assign T2374 = $signed(30'h11f56d44) * $signed(16'h0);
  assign T2375 = T2373[6'h2d:6'h2d];
  assign T2376 = $signed(T2377) / $signed(22'h100000);
  assign T2377 = $signed(31'h3d6dbf43) * $signed(16'h1);
  assign T2378 = T1637[1'h0:1'h0];
  assign T2379 = T1637[1'h1:1'h1];
  assign T2380 = T2409 ? T2395 : T2381;
  assign T2381 = T2394 ? twiddle3_1_13_real : twiddle3_1_12_real;
  assign twiddle3_1_12_real = T2386 + T2382;
  assign T2382 = {T2385, T2383};
  assign T2383 = $signed(T2384) / $signed(22'h100000);
  assign T2384 = $signed(30'h138a760d) * $signed(16'h0);
  assign T2385 = T2383[6'h2d:6'h2d];
  assign T2386 = $signed(T2387) / $signed(22'h100000);
  assign T2387 = $signed(31'h3cf1a11d) * $signed(16'h1);
  assign twiddle3_1_13_real = T2392 + T2388;
  assign T2388 = {T2391, T2389};
  assign T2389 = $signed(T2390) / $signed(22'h100000);
  assign T2390 = $signed(30'h151c26b1) * $signed(16'h0);
  assign T2391 = T2389[6'h2d:6'h2d];
  assign T2392 = $signed(T2393) / $signed(22'h100000);
  assign T2393 = $signed(31'h3c6b14d5) * $signed(16'h1);
  assign T2394 = T1637[1'h0:1'h0];
  assign T2395 = T2408 ? twiddle3_1_15_real : twiddle3_1_14_real;
  assign twiddle3_1_14_real = T2400 + T2396;
  assign T2396 = {T2399, T2397};
  assign T2397 = $signed(T2398) / $signed(22'h100000);
  assign T2398 = $signed(30'h16aa3a72) * $signed(16'h0);
  assign T2399 = T2397[6'h2d:6'h2d];
  assign T2400 = $signed(T2401) / $signed(22'h100000);
  assign T2401 = $signed(31'h3bda3171) * $signed(16'h1);
  assign twiddle3_1_15_real = T2406 + T2402;
  assign T2402 = {T2405, T2403};
  assign T2403 = $signed(T2404) / $signed(22'h100000);
  assign T2404 = $signed(30'h18346d2d) * $signed(16'h0);
  assign T2405 = T2403[6'h2d:6'h2d];
  assign T2406 = $signed(T2407) / $signed(22'h100000);
  assign T2407 = $signed(31'h3b3f0fbf) * $signed(16'h1);
  assign T2408 = T1637[1'h0:1'h0];
  assign T2409 = T1637[1'h1:1'h1];
  assign T2410 = T1637[2'h2:2'h2];
  assign T2411 = T2347[6'h2e:6'h2e];
  assign T2412 = T1637[2'h3:2'h3];
  assign T2413 = {T2518, T2414};
  assign T2414 = T2517 ? T2471 : T2415;
  assign T2415 = T2470 ? T2446 : T2416;
  assign T2416 = T2445 ? T2431 : T2417;
  assign T2417 = T2430 ? twiddle3_1_17_real : twiddle3_1_16_real;
  assign twiddle3_1_16_real = T2422 + T2418;
  assign T2418 = {T2421, T2419};
  assign T2419 = $signed(T2420) / $signed(22'h100000);
  assign T2420 = $signed(30'h19ba7b6c) * $signed(16'h0);
  assign T2421 = T2419[6'h2d:6'h2d];
  assign T2422 = $signed(T2423) / $signed(22'h100000);
  assign T2423 = $signed(31'h3a99ca4a) * $signed(16'h1);
  assign twiddle3_1_17_real = T2428 + T2424;
  assign T2424 = {T2427, T2425};
  assign T2425 = $signed(T2426) / $signed(22'h100000);
  assign T2426 = $signed(30'h1b3c226e) * $signed(16'h0);
  assign T2427 = T2425[6'h2d:6'h2d];
  assign T2428 = $signed(T2429) / $signed(22'h100000);
  assign T2429 = $signed(31'h39ea7d5c) * $signed(16'h1);
  assign T2430 = T1637[1'h0:1'h0];
  assign T2431 = T2444 ? twiddle3_1_19_real : twiddle3_1_18_real;
  assign twiddle3_1_18_real = T2436 + T2432;
  assign T2432 = {T2435, T2433};
  assign T2433 = $signed(T2434) / $signed(22'h100000);
  assign T2434 = $signed(30'h1cb92032) * $signed(16'h0);
  assign T2435 = T2433[6'h2d:6'h2d];
  assign T2436 = $signed(T2437) / $signed(22'h100000);
  assign T2437 = $signed(31'h393146f5) * $signed(16'h1);
  assign twiddle3_1_19_real = T2442 + T2438;
  assign T2438 = {T2441, T2439};
  assign T2439 = $signed(T2440) / $signed(22'h100000);
  assign T2440 = $signed(30'h1e313383) * $signed(16'h0);
  assign T2441 = T2439[6'h2d:6'h2d];
  assign T2442 = $signed(T2443) / $signed(22'h100000);
  assign T2443 = $signed(31'h386e46c7) * $signed(16'h1);
  assign T2444 = T1637[1'h0:1'h0];
  assign T2445 = T1637[1'h1:1'h1];
  assign T2446 = T2469 ? T2459 : T2447;
  assign T2447 = T2458 ? twiddle3_1_21_real : twiddle3_1_20_real;
  assign twiddle3_1_20_real = T2452 + T2448;
  assign T2448 = {T2451, T2449};
  assign T2449 = $signed(T2450) / $signed(22'h100000);
  assign T2450 = $signed(30'h1fa41c05) * $signed(16'h0);
  assign T2451 = T2449[6'h2d:6'h2d];
  assign T2452 = $signed(T2453) / $signed(22'h100000);
  assign T2453 = $signed(31'h37a19e34) * $signed(16'h1);
  assign twiddle3_1_21_real = T2456 + T2454;
  assign T2454 = $signed(T2455) / $signed(22'h100000);
  assign T2455 = $signed(31'h21119a3d) * $signed(16'h0);
  assign T2456 = $signed(T2457) / $signed(22'h100000);
  assign T2457 = $signed(31'h36cb7040) * $signed(16'h1);
  assign T2458 = T1637[1'h0:1'h0];
  assign T2459 = T2468 ? twiddle3_1_23_real : twiddle3_1_22_real;
  assign twiddle3_1_22_real = T2462 + T2460;
  assign T2460 = $signed(T2461) / $signed(22'h100000);
  assign T2461 = $signed(31'h22796f9d) * $signed(16'h0);
  assign T2462 = $signed(T2463) / $signed(22'h100000);
  assign T2463 = $signed(31'h35ebe194) * $signed(16'h1);
  assign twiddle3_1_23_real = T2466 + T2464;
  assign T2464 = $signed(T2465) / $signed(22'h100000);
  assign T2465 = $signed(31'h23db5e91) * $signed(16'h0);
  assign T2466 = $signed(T2467) / $signed(22'h100000);
  assign T2467 = $signed(31'h35031873) * $signed(16'h1);
  assign T2468 = T1637[1'h0:1'h0];
  assign T2469 = T1637[1'h1:1'h1];
  assign T2470 = T1637[2'h2:2'h2];
  assign T2471 = T2516 ? T2494 : T2472;
  assign T2472 = T2493 ? T2483 : T2473;
  assign T2473 = T2482 ? twiddle3_1_25_real : twiddle3_1_24_real;
  assign twiddle3_1_24_real = T2476 + T2474;
  assign T2474 = $signed(T2475) / $signed(22'h100000);
  assign T2475 = $signed(31'h25372a85) * $signed(16'h0);
  assign T2476 = $signed(T2477) / $signed(22'h100000);
  assign T2477 = $signed(31'h34113cb3) * $signed(16'h1);
  assign twiddle3_1_25_real = T2480 + T2478;
  assign T2478 = $signed(T2479) / $signed(22'h100000);
  assign T2479 = $signed(31'h268c97f3) * $signed(16'h0);
  assign T2480 = $signed(T2481) / $signed(22'h100000);
  assign T2481 = $signed(31'h331677ba) * $signed(16'h1);
  assign T2482 = T1637[1'h0:1'h0];
  assign T2483 = T2492 ? twiddle3_1_27_real : twiddle3_1_26_real;
  assign twiddle3_1_26_real = T2486 + T2484;
  assign T2484 = $signed(T2485) / $signed(22'h100000);
  assign T2485 = $signed(31'h27db6c6d) * $signed(16'h0);
  assign T2486 = $signed(T2487) / $signed(22'h100000);
  assign T2487 = $signed(31'h3212f472) * $signed(16'h1);
  assign twiddle3_1_27_real = T2490 + T2488;
  assign T2488 = $signed(T2489) / $signed(22'h100000);
  assign T2489 = $signed(31'h29236ea4) * $signed(16'h0);
  assign T2490 = $signed(T2491) / $signed(22'h100000);
  assign T2491 = $signed(31'h3106df45) * $signed(16'h1);
  assign T2492 = T1637[1'h0:1'h0];
  assign T2493 = T1637[1'h1:1'h1];
  assign T2494 = T2515 ? T2505 : T2495;
  assign T2495 = T2504 ? twiddle3_1_29_real : twiddle3_1_28_real;
  assign twiddle3_1_28_real = T2498 + T2496;
  assign T2496 = $signed(T2497) / $signed(22'h100000);
  assign T2497 = $signed(31'h2a646676) * $signed(16'h0);
  assign T2498 = $signed(T2499) / $signed(22'h100000);
  assign T2499 = $signed(31'h2ff26615) * $signed(16'h1);
  assign twiddle3_1_29_real = T2502 + T2500;
  assign T2500 = $signed(T2501) / $signed(22'h100000);
  assign T2501 = $signed(31'h2b9e1cf3) * $signed(16'h0);
  assign T2502 = $signed(T2503) / $signed(22'h100000);
  assign T2503 = $signed(31'h2ed5b833) * $signed(16'h1);
  assign T2504 = T1637[1'h0:1'h0];
  assign T2505 = T2514 ? twiddle3_1_31_real : twiddle3_1_30_real;
  assign twiddle3_1_30_real = T2508 + T2506;
  assign T2506 = $signed(T2507) / $signed(22'h100000);
  assign T2507 = $signed(31'h2cd05c6c) * $signed(16'h0);
  assign T2508 = $signed(T2509) / $signed(22'h100000);
  assign T2509 = $signed(31'h2db10657) * $signed(16'h1);
  assign twiddle3_1_31_real = T2512 + T2510;
  assign T2510 = $signed(T2511) / $signed(22'h100000);
  assign T2511 = $signed(31'h2dfaf076) * $signed(16'h0);
  assign T2512 = $signed(T2513) / $signed(22'h100000);
  assign T2513 = $signed(31'h2c848299) * $signed(16'h1);
  assign T2514 = T1637[1'h0:1'h0];
  assign T2515 = T1637[1'h1:1'h1];
  assign T2516 = T1637[2'h2:2'h2];
  assign T2517 = T1637[2'h3:2'h3];
  assign T2518 = T2414[6'h2e:6'h2e];
  assign T2519 = T1637[3'h4:3'h4];
  assign T2520 = {T2770, T2521};
  assign T2521 = T2769 ? T2630 : T2522;
  assign T2522 = T2629 ? T2569 : T2523;
  assign T2523 = T2568 ? T2546 : T2524;
  assign T2524 = T2545 ? T2535 : T2525;
  assign T2525 = T2534 ? twiddle3_1_33_real : twiddle3_1_32_real;
  assign twiddle3_1_32_real = T2528 + T2526;
  assign T2526 = $signed(T2527) / $signed(22'h100000);
  assign T2527 = $signed(31'h2f1da5f8) * $signed(16'h0);
  assign T2528 = $signed(T2529) / $signed(22'h100000);
  assign T2529 = $signed(31'h2b506069) * $signed(16'h1);
  assign twiddle3_1_33_real = T2532 + T2530;
  assign T2530 = $signed(T2531) / $signed(22'h100000);
  assign T2531 = $signed(31'h30384b31) * $signed(16'h0);
  assign T2532 = $signed(T2533) / $signed(22'h100000);
  assign T2533 = $signed(31'h2a14d481) * $signed(16'h1);
  assign T2534 = T1637[1'h0:1'h0];
  assign T2535 = T2544 ? twiddle3_1_35_real : twiddle3_1_34_real;
  assign twiddle3_1_34_real = T2538 + T2536;
  assign T2536 = $signed(T2537) / $signed(22'h100000);
  assign T2537 = $signed(31'h314aafc2) * $signed(16'h0);
  assign T2538 = $signed(T2539) / $signed(22'h100000);
  assign T2539 = $signed(31'h28d214e4) * $signed(16'h1);
  assign twiddle3_1_35_real = T2542 + T2540;
  assign T2540 = $signed(T2541) / $signed(22'h100000);
  assign T2541 = $signed(31'h3254a4b4) * $signed(16'h0);
  assign T2542 = $signed(T2543) / $signed(22'h100000);
  assign T2543 = $signed(31'h278858cd) * $signed(16'h1);
  assign T2544 = T1637[1'h0:1'h0];
  assign T2545 = T1637[1'h1:1'h1];
  assign T2546 = T2567 ? T2557 : T2547;
  assign T2547 = T2556 ? twiddle3_1_37_real : twiddle3_1_36_real;
  assign twiddle3_1_36_real = T2550 + T2548;
  assign T2548 = $signed(T2549) / $signed(22'h100000);
  assign T2549 = $signed(31'h3355fc84) * $signed(16'h0);
  assign T2550 = $signed(T2551) / $signed(22'h100000);
  assign T2551 = $signed(31'h2637d8ab) * $signed(16'h1);
  assign twiddle3_1_37_real = T2554 + T2552;
  assign T2552 = $signed(T2553) / $signed(22'h100000);
  assign T2553 = $signed(31'h344e8b25) * $signed(16'h0);
  assign T2554 = $signed(T2555) / $signed(22'h100000);
  assign T2555 = $signed(31'h24e0ce16) * $signed(16'h1);
  assign T2556 = T1637[1'h0:1'h0];
  assign T2557 = T2566 ? twiddle3_1_39_real : twiddle3_1_38_real;
  assign twiddle3_1_38_real = T2560 + T2558;
  assign T2558 = $signed(T2559) / $signed(22'h100000);
  assign T2559 = $signed(31'h353e260f) * $signed(16'h0);
  assign T2560 = $signed(T2561) / $signed(22'h100000);
  assign T2561 = $signed(31'h238373c3) * $signed(16'h1);
  assign twiddle3_1_39_real = T2564 + T2562;
  assign T2562 = $signed(T2563) / $signed(22'h100000);
  assign T2563 = $signed(31'h3624a440) * $signed(16'h0);
  assign T2564 = $signed(T2565) / $signed(22'h100000);
  assign T2565 = $signed(31'h2220057c) * $signed(16'h1);
  assign T2566 = T1637[1'h0:1'h0];
  assign T2567 = T1637[1'h1:1'h1];
  assign T2568 = T1637[2'h2:2'h2];
  assign T2569 = T2628 ? T2598 : T2570;
  assign T2570 = T2597 ? T2583 : T2571;
  assign T2571 = T2582 ? twiddle3_1_41_real : twiddle3_1_40_real;
  assign twiddle3_1_40_real = T2574 + T2572;
  assign T2572 = $signed(T2573) / $signed(22'h100000);
  assign T2573 = $signed(31'h3701de44) * $signed(16'h0);
  assign T2574 = $signed(T2575) / $signed(22'h100000);
  assign T2575 = $signed(31'h20b6c016) * $signed(16'h1);
  assign twiddle3_1_41_real = T2578 + T2576;
  assign T2576 = $signed(T2577) / $signed(22'h100000);
  assign T2577 = $signed(31'h37d5ae3f) * $signed(16'h0);
  assign T2578 = {T2581, T2579};
  assign T2579 = $signed(T2580) / $signed(22'h100000);
  assign T2580 = $signed(30'h1f47e165) * $signed(16'h1);
  assign T2581 = T2579[6'h2d:6'h2d];
  assign T2582 = T1637[1'h0:1'h0];
  assign T2583 = T2596 ? twiddle3_1_43_real : twiddle3_1_42_real;
  assign twiddle3_1_42_real = T2586 + T2584;
  assign T2584 = $signed(T2585) / $signed(22'h100000);
  assign T2585 = $signed(31'h389feff1) * $signed(16'h0);
  assign T2586 = {T2589, T2587};
  assign T2587 = $signed(T2588) / $signed(22'h100000);
  assign T2588 = $signed(30'h1dd3a832) * $signed(16'h1);
  assign T2589 = T2587[6'h2d:6'h2d];
  assign twiddle3_1_43_real = T2592 + T2590;
  assign T2590 = $signed(T2591) / $signed(22'h100000);
  assign T2591 = $signed(31'h396080bd) * $signed(16'h0);
  assign T2592 = {T2595, T2593};
  assign T2593 = $signed(T2594) / $signed(22'h100000);
  assign T2594 = $signed(30'h1c5a5433) * $signed(16'h1);
  assign T2595 = T2593[6'h2d:6'h2d];
  assign T2596 = T1637[1'h0:1'h0];
  assign T2597 = T1637[1'h1:1'h1];
  assign T2598 = T2627 ? T2613 : T2599;
  assign T2599 = T2612 ? twiddle3_1_45_real : twiddle3_1_44_real;
  assign twiddle3_1_44_real = T2602 + T2600;
  assign T2600 = $signed(T2601) / $signed(22'h100000);
  assign T2601 = $signed(31'h3a173fae) * $signed(16'h0);
  assign T2602 = {T2605, T2603};
  assign T2603 = $signed(T2604) / $signed(22'h100000);
  assign T2604 = $signed(30'h1adc25fb) * $signed(16'h1);
  assign T2605 = T2603[6'h2d:6'h2d];
  assign twiddle3_1_45_real = T2608 + T2606;
  assign T2606 = $signed(T2607) / $signed(22'h100000);
  assign T2607 = $signed(31'h3ac40d7d) * $signed(16'h0);
  assign T2608 = {T2611, T2609};
  assign T2609 = $signed(T2610) / $signed(22'h100000);
  assign T2610 = $signed(30'h19595ef2) * $signed(16'h1);
  assign T2611 = T2609[6'h2d:6'h2d];
  assign T2612 = T1637[1'h0:1'h0];
  assign T2613 = T2626 ? twiddle3_1_47_real : twiddle3_1_46_real;
  assign twiddle3_1_46_real = T2616 + T2614;
  assign T2614 = $signed(T2615) / $signed(22'h100000);
  assign T2615 = $signed(31'h3b66cc97) * $signed(16'h0);
  assign T2616 = {T2619, T2617};
  assign T2617 = $signed(T2618) / $signed(22'h100000);
  assign T2618 = $signed(30'h17d2414a) * $signed(16'h1);
  assign T2619 = T2617[6'h2d:6'h2d];
  assign twiddle3_1_47_real = T2622 + T2620;
  assign T2620 = $signed(T2621) / $signed(22'h100000);
  assign T2621 = $signed(31'h3bff6121) * $signed(16'h0);
  assign T2622 = {T2625, T2623};
  assign T2623 = $signed(T2624) / $signed(22'h100000);
  assign T2624 = $signed(30'h16470ff4) * $signed(16'h1);
  assign T2625 = T2623[6'h2d:6'h2d];
  assign T2626 = T1637[1'h0:1'h0];
  assign T2627 = T1637[1'h1:1'h1];
  assign T2628 = T1637[2'h2:2'h2];
  assign T2629 = T1637[2'h3:2'h3];
  assign T2630 = T2768 ? T2698 : T2631;
  assign T2631 = T2697 ? T2663 : T2632;
  assign T2632 = T2662 ? T2647 : T2633;
  assign T2633 = T2646 ? twiddle3_1_49_real : twiddle3_1_48_real;
  assign twiddle3_1_48_real = T2636 + T2634;
  assign T2634 = $signed(T2635) / $signed(22'h100000);
  assign T2635 = $signed(31'h3c8db0ff) * $signed(16'h0);
  assign T2636 = {T2639, T2637};
  assign T2637 = $signed(T2638) / $signed(22'h100000);
  assign T2638 = $signed(30'h14b80e91) * $signed(16'h1);
  assign T2639 = T2637[6'h2d:6'h2d];
  assign twiddle3_1_49_real = T2642 + T2640;
  assign T2640 = $signed(T2641) / $signed(22'h100000);
  assign T2641 = $signed(31'h3d11a3d6) * $signed(16'h0);
  assign T2642 = {T2645, T2643};
  assign T2643 = $signed(T2644) / $signed(22'h100000);
  assign T2644 = $signed(30'h1325816c) * $signed(16'h1);
  assign T2645 = T2643[6'h2d:6'h2d];
  assign T2646 = T1637[1'h0:1'h0];
  assign T2647 = T2661 ? twiddle3_1_51_real : twiddle3_1_50_real;
  assign twiddle3_1_50_real = T2650 + T2648;
  assign T2648 = $signed(T2649) / $signed(22'h100000);
  assign T2649 = $signed(31'h3d8b2310) * $signed(16'h0);
  assign T2650 = {T2653, T2651};
  assign T2651 = $signed(T2652) / $signed(22'h100000);
  assign T2652 = $signed(30'h118fad69) * $signed(16'h1);
  assign T2653 = T2651[6'h2d:6'h2d];
  assign twiddle3_1_51_real = T2656 + T2654;
  assign T2654 = $signed(T2655) / $signed(22'h100000);
  assign T2655 = $signed(31'h3dfa19e2) * $signed(16'h0);
  assign T2656 = {T2659, T2657};
  assign T2657 = $signed(T2658) / $signed(22'h100000);
  assign T2658 = $signed(29'hff6d7fd) * $signed(16'h1);
  assign T2659 = T2660 ? 2'h3 : 2'h0;
  assign T2660 = T2657[6'h2c:6'h2c];
  assign T2661 = T1637[1'h0:1'h0];
  assign T2662 = T1637[1'h1:1'h1];
  assign T2663 = T2696 ? T2680 : T2664;
  assign T2664 = T2679 ? twiddle3_1_53_real : twiddle3_1_52_real;
  assign twiddle3_1_52_real = T2667 + T2665;
  assign T2665 = $signed(T2666) / $signed(22'h100000);
  assign T2666 = $signed(31'h3e5e754f) * $signed(16'h0);
  assign T2667 = {T2670, T2668};
  assign T2668 = $signed(T2669) / $signed(22'h100000);
  assign T2669 = $signed(29'he5b4720) * $signed(16'h1);
  assign T2670 = T2671 ? 2'h3 : 2'h0;
  assign T2671 = T2668[6'h2c:6'h2c];
  assign twiddle3_1_53_real = T2674 + T2672;
  assign T2672 = $signed(T2673) / $signed(22'h100000);
  assign T2673 = $signed(31'h3eb8242a) * $signed(16'h0);
  assign T2674 = {T2677, T2675};
  assign T2675 = $signed(T2676) / $signed(22'h100000);
  assign T2676 = $signed(29'hcbd4142) * $signed(16'h1);
  assign T2677 = T2678 ? 2'h3 : 2'h0;
  assign T2678 = T2675[6'h2c:6'h2c];
  assign T2679 = T1637[1'h0:1'h0];
  assign T2680 = T2695 ? twiddle3_1_55_real : twiddle3_1_54_real;
  assign twiddle3_1_54_real = T2683 + T2681;
  assign T2681 = $signed(T2682) / $signed(22'h100000);
  assign T2682 = $signed(31'h3f071719) * $signed(16'h0);
  assign T2683 = {T2686, T2684};
  assign T2684 = $signed(T2685) / $signed(22'h100000);
  assign T2685 = $signed(29'hb1d0d3f) * $signed(16'h1);
  assign T2686 = T2687 ? 2'h3 : 2'h0;
  assign T2687 = T2684[6'h2c:6'h2c];
  assign twiddle3_1_55_real = T2690 + T2688;
  assign T2688 = $signed(T2689) / $signed(22'h100000);
  assign T2689 = $signed(31'h3f4b4099) * $signed(16'h0);
  assign T2690 = {T2693, T2691};
  assign T2691 = $signed(T2692) / $signed(22'h100000);
  assign T2692 = $signed(29'h97af251) * $signed(16'h1);
  assign T2693 = T2694 ? 2'h3 : 2'h0;
  assign T2694 = T2691[6'h2c:6'h2c];
  assign T2695 = T1637[1'h0:1'h0];
  assign T2696 = T1637[1'h1:1'h1];
  assign T2697 = T1637[2'h2:2'h2];
  assign T2698 = T2767 ? T2733 : T2699;
  assign T2699 = T2732 ? T2716 : T2700;
  assign T2700 = T2715 ? twiddle3_1_57_real : twiddle3_1_56_real;
  assign twiddle3_1_56_real = T2703 + T2701;
  assign T2701 = $signed(T2702) / $signed(22'h100000);
  assign T2702 = $signed(31'h3f849500) * $signed(16'h0);
  assign T2703 = {T2706, T2704};
  assign T2704 = $signed(T2705) / $signed(22'h100000);
  assign T2705 = $signed(28'h7d73808) * $signed(16'h1);
  assign T2706 = T2707 ? 3'h7 : 3'h0;
  assign T2707 = T2704[6'h2b:6'h2b];
  assign twiddle3_1_57_real = T2710 + T2708;
  assign T2708 = $signed(T2709) / $signed(22'h100000);
  assign T2709 = $signed(31'h3fb30a7f) * $signed(16'h0);
  assign T2710 = {T2713, T2711};
  assign T2711 = $signed(T2712) / $signed(22'h100000);
  assign T2712 = $signed(28'h6322638) * $signed(16'h1);
  assign T2713 = T2714 ? 3'h7 : 3'h0;
  assign T2714 = T2711[6'h2b:6'h2b];
  assign T2715 = T1637[1'h0:1'h0];
  assign T2716 = T2731 ? twiddle3_1_59_real : twiddle3_1_58_real;
  assign twiddle3_1_58_real = T2719 + T2717;
  assign T2717 = $signed(T2718) / $signed(22'h100000);
  assign T2718 = $signed(31'h3fd69921) * $signed(16'h0);
  assign T2719 = {T2722, T2720};
  assign T2720 = $signed(T2721) / $signed(22'h100000);
  assign T2721 = $signed(28'h48c04f3) * $signed(16'h1);
  assign T2722 = T2723 ? 3'h7 : 3'h0;
  assign T2723 = T2720[6'h2b:6'h2b];
  assign twiddle3_1_59_real = T2726 + T2724;
  assign T2724 = $signed(T2725) / $signed(22'h100000);
  assign T2725 = $signed(31'h3fef3ad1) * $signed(16'h0);
  assign T2726 = {T2729, T2727};
  assign T2727 = $signed(T2728) / $signed(22'h100000);
  assign T2728 = $signed(27'h2e51c76) * $signed(16'h1);
  assign T2729 = T2730 ? 4'hf : 4'h0;
  assign T2730 = T2727[6'h2a:6'h2a];
  assign T2731 = T1637[1'h0:1'h0];
  assign T2732 = T1637[1'h1:1'h1];
  assign T2733 = T2766 ? T2750 : T2734;
  assign T2734 = T2749 ? twiddle3_1_61_real : twiddle3_1_60_real;
  assign twiddle3_1_60_real = T2737 + T2735;
  assign T2735 = $signed(T2736) / $signed(22'h100000);
  assign T2736 = $signed(31'h3ffceb58) * $signed(16'h0);
  assign T2737 = {T2740, T2738};
  assign T2738 = $signed(T2739) / $signed(22'h100000);
  assign T2739 = $signed(26'h13db523) * $signed(16'h1);
  assign T2740 = T2741 ? 5'h1f : 5'h0;
  assign T2741 = T2738[6'h29:6'h29];
  assign twiddle3_1_61_real = T2744 + T2742;
  assign T2742 = $signed(T2743) / $signed(22'h100000);
  assign T2743 = $signed(31'h3fffa85e) * $signed(16'h0);
  assign T2744 = {T2747, T2745};
  assign T2745 = $signed(T2746) / $signed(22'h100000);
  assign T2746 = $signed(24'h961772) * $signed(16'h1);
  assign T2747 = T2748 ? 7'h7f : 7'h0;
  assign T2748 = T2745[6'h27:6'h27];
  assign T2749 = T1637[1'h0:1'h0];
  assign T2750 = T2765 ? twiddle3_1_63_real : twiddle3_1_62_real;
  assign twiddle3_1_62_real = T2753 + T2751;
  assign T2751 = $signed(T2752) / $signed(22'h100000);
  assign T2752 = $signed(31'h3ff7716b) * $signed(16'h0);
  assign T2753 = {T2756, T2754};
  assign T2754 = $signed(T2755) / $signed(22'h100000);
  assign T2755 = $signed(27'h5ee8bdf) * $signed(16'h1);
  assign T2756 = T2757 ? 4'hf : 4'h0;
  assign T2757 = T2754[6'h2a:6'h2a];
  assign twiddle3_1_63_real = T2760 + T2758;
  assign T2758 = $signed(T2759) / $signed(22'h100000);
  assign T2759 = $signed(31'h3fe447e6) * $signed(16'h0);
  assign T2760 = {T2763, T2761};
  assign T2761 = $signed(T2762) / $signed(22'h100000);
  assign T2762 = $signed(27'h4475aea) * $signed(16'h1);
  assign T2763 = T2764 ? 4'hf : 4'h0;
  assign T2764 = T2761[6'h2a:6'h2a];
  assign T2765 = T1637[1'h0:1'h0];
  assign T2766 = T1637[1'h1:1'h1];
  assign T2767 = T1637[2'h2:2'h2];
  assign T2768 = T1637[2'h3:2'h3];
  assign T2769 = T1637[3'h4:3'h4];
  assign T2770 = T2521[6'h2e:6'h2e];
  assign T2771 = T1637[3'h5:3'h5];
  assign T2772 = {T2914, T2773};
  assign T2773 = T2913 ? twiddle3_1_80_real : T2774;
  assign T2774 = T2906 ? T2844 : T2775;
  assign T2775 = T2843 ? T2810 : T2776;
  assign T2776 = T2809 ? T2793 : T2777;
  assign T2777 = T2792 ? twiddle3_1_65_real : twiddle3_1_64_real;
  assign twiddle3_1_64_real = T2780 + T2778;
  assign T2778 = $signed(T2779) / $signed(22'h100000);
  assign T2779 = $signed(31'h3fc62f18) * $signed(16'h0);
  assign T2780 = {T2783, T2781};
  assign T2781 = $signed(T2782) / $signed(22'h100000);
  assign T2782 = $signed(28'haa0ccff) * $signed(16'h1);
  assign T2783 = T2784 ? 3'h7 : 3'h0;
  assign T2784 = T2781[6'h2b:6'h2b];
  assign twiddle3_1_65_real = T2787 + T2785;
  assign T2785 = $signed(T2786) / $signed(22'h100000);
  assign T2786 = $signed(31'h3f9d2c27) * $signed(16'h0);
  assign T2787 = {T2790, T2788};
  assign T2788 = $signed(T2789) / $signed(22'h100000);
  assign T2789 = $signed(28'h8fb2a6f) * $signed(16'h1);
  assign T2790 = T2791 ? 3'h7 : 3'h0;
  assign T2791 = T2788[6'h2b:6'h2b];
  assign T2792 = T1637[1'h0:1'h0];
  assign T2793 = T2808 ? twiddle3_1_67_real : twiddle3_1_66_real;
  assign twiddle3_1_66_real = T2796 + T2794;
  assign T2794 = $signed(T2795) / $signed(22'h100000);
  assign T2795 = $signed(31'h3f694618) * $signed(16'h0);
  assign T2796 = {T2799, T2797};
  assign T2797 = $signed(T2798) / $signed(22'h100000);
  assign T2798 = $signed(29'h1756bb64) * $signed(16'h1);
  assign T2799 = T2800 ? 2'h3 : 2'h0;
  assign T2800 = T2797[6'h2c:6'h2c];
  assign twiddle3_1_67_real = T2803 + T2801;
  assign T2801 = $signed(T2802) / $signed(22'h100000);
  assign T2802 = $signed(31'h3f2a85cc) * $signed(16'h0);
  assign T2803 = {T2806, T2804};
  assign T2804 = $signed(T2805) / $signed(22'h100000);
  assign T2805 = $signed(29'h15b3c7d2) * $signed(16'h1);
  assign T2806 = T2807 ? 2'h3 : 2'h0;
  assign T2807 = T2804[6'h2c:6'h2c];
  assign T2808 = T1637[1'h0:1'h0];
  assign T2809 = T1637[1'h1:1'h1];
  assign T2810 = T2842 ? T2827 : T2811;
  assign T2811 = T2826 ? twiddle3_1_69_real : twiddle3_1_68_real;
  assign twiddle3_1_68_real = T2814 + T2812;
  assign T2812 = $signed(T2813) / $signed(22'h100000);
  assign T2813 = $signed(31'h3ee0f602) * $signed(16'h0);
  assign T2814 = {T2817, T2815};
  assign T2815 = $signed(T2816) / $signed(22'h100000);
  assign T2816 = $signed(29'h1412976d) * $signed(16'h1);
  assign T2817 = T2818 ? 2'h3 : 2'h0;
  assign T2818 = T2815[6'h2c:6'h2c];
  assign twiddle3_1_69_real = T2821 + T2819;
  assign T2819 = $signed(T2820) / $signed(22'h100000);
  assign T2820 = $signed(31'h3e8ca34f) * $signed(16'h0);
  assign T2821 = {T2824, T2822};
  assign T2822 = $signed(T2823) / $signed(22'h100000);
  assign T2823 = $signed(29'h1273719b) * $signed(16'h1);
  assign T2824 = T2825 ? 2'h3 : 2'h0;
  assign T2825 = T2822[6'h2c:6'h2c];
  assign T2826 = T1637[1'h0:1'h0];
  assign T2827 = T2841 ? twiddle3_1_71_real : twiddle3_1_70_real;
  assign twiddle3_1_70_real = T2830 + T2828;
  assign T2828 = $signed(T2829) / $signed(22'h100000);
  assign T2829 = $signed(31'h3e2d9c23) * $signed(16'h0);
  assign T2830 = {T2833, T2831};
  assign T2831 = $signed(T2832) / $signed(22'h100000);
  assign T2832 = $signed(29'h10d69d68) * $signed(16'h1);
  assign T2833 = T2834 ? 2'h3 : 2'h0;
  assign T2834 = T2831[6'h2c:6'h2c];
  assign twiddle3_1_71_real = T2837 + T2835;
  assign T2835 = $signed(T2836) / $signed(22'h100000);
  assign T2836 = $signed(31'h3dc3f0c1) * $signed(16'h0);
  assign T2837 = {T2840, T2838};
  assign T2838 = $signed(T2839) / $signed(22'h100000);
  assign T2839 = $signed(30'h2f3c617d) * $signed(16'h1);
  assign T2840 = T2838[6'h2d:6'h2d];
  assign T2841 = T1637[1'h0:1'h0];
  assign T2842 = T1637[1'h1:1'h1];
  assign T2843 = T1637[2'h2:2'h2];
  assign T2844 = T2905 ? T2875 : T2845;
  assign T2845 = T2874 ? T2860 : T2846;
  assign T2846 = T2859 ? twiddle3_1_73_real : twiddle3_1_72_real;
  assign twiddle3_1_72_real = T2849 + T2847;
  assign T2847 = $signed(T2848) / $signed(22'h100000);
  assign T2848 = $signed(31'h3d4fb33e) * $signed(16'h0);
  assign T2849 = {T2852, T2850};
  assign T2850 = $signed(T2851) / $signed(22'h100000);
  assign T2851 = $signed(30'h2da5040e) * $signed(16'h1);
  assign T2852 = T2850[6'h2d:6'h2d];
  assign twiddle3_1_73_real = T2855 + T2853;
  assign T2853 = $signed(T2854) / $signed(22'h100000);
  assign T2854 = $signed(31'h3cd0f77f) * $signed(16'h0);
  assign T2855 = {T2858, T2856};
  assign T2856 = $signed(T2857) / $signed(22'h100000);
  assign T2857 = $signed(30'h2c10cad4) * $signed(16'h1);
  assign T2858 = T2856[6'h2d:6'h2d];
  assign T2859 = T1637[1'h0:1'h0];
  assign T2860 = T2873 ? twiddle3_1_75_real : twiddle3_1_74_real;
  assign twiddle3_1_74_real = T2863 + T2861;
  assign T2861 = $signed(T2862) / $signed(22'h100000);
  assign T2862 = $signed(31'h3c47d336) * $signed(16'h0);
  assign T2863 = {T2866, T2864};
  assign T2864 = $signed(T2865) / $signed(22'h100000);
  assign T2865 = $signed(30'h2a7ffafd) * $signed(16'h1);
  assign T2866 = T2864[6'h2d:6'h2d];
  assign twiddle3_1_75_real = T2869 + T2867;
  assign T2867 = $signed(T2868) / $signed(22'h100000);
  assign T2868 = $signed(31'h3bb45dda) * $signed(16'h0);
  assign T2869 = {T2872, T2870};
  assign T2870 = $signed(T2871) / $signed(22'h100000);
  assign T2871 = $signed(30'h28f2d921) * $signed(16'h1);
  assign T2872 = T2870[6'h2d:6'h2d];
  assign T2873 = T1637[1'h0:1'h0];
  assign T2874 = T1637[1'h1:1'h1];
  assign T2875 = T2904 ? T2890 : T2876;
  assign T2876 = T2889 ? twiddle3_1_77_real : twiddle3_1_76_real;
  assign twiddle3_1_76_real = T2879 + T2877;
  assign T2877 = $signed(T2878) / $signed(22'h100000);
  assign T2878 = $signed(31'h3b16b0a8) * $signed(16'h0);
  assign T2879 = {T2882, T2880};
  assign T2880 = $signed(T2881) / $signed(22'h100000);
  assign T2881 = $signed(30'h2769a939) * $signed(16'h1);
  assign T2882 = T2880[6'h2d:6'h2d];
  assign twiddle3_1_77_real = T2885 + T2883;
  assign T2883 = $signed(T2884) / $signed(22'h100000);
  assign T2884 = $signed(31'h3a6ee69d) * $signed(16'h0);
  assign T2885 = {T2888, T2886};
  assign T2886 = $signed(T2887) / $signed(22'h100000);
  assign T2887 = $signed(30'h25e4ae8e) * $signed(16'h1);
  assign T2888 = T2886[6'h2d:6'h2d];
  assign T2889 = T1637[1'h0:1'h0];
  assign T2890 = T2903 ? twiddle3_1_79_real : twiddle3_1_78_real;
  assign twiddle3_1_78_real = T2893 + T2891;
  assign T2891 = $signed(T2892) / $signed(22'h100000);
  assign T2892 = $signed(31'h39bd1c70) * $signed(16'h0);
  assign T2893 = {T2896, T2894};
  assign T2894 = $signed(T2895) / $signed(22'h100000);
  assign T2895 = $signed(30'h24642bb3) * $signed(16'h1);
  assign T2896 = T2894[6'h2d:6'h2d];
  assign twiddle3_1_79_real = T2899 + T2897;
  assign T2897 = $signed(T2898) / $signed(22'h100000);
  assign T2898 = $signed(31'h3901708e) * $signed(16'h0);
  assign T2899 = {T2902, T2900};
  assign T2900 = $signed(T2901) / $signed(22'h100000);
  assign T2901 = $signed(30'h22e86278) * $signed(16'h1);
  assign T2902 = T2900[6'h2d:6'h2d];
  assign T2903 = T1637[1'h0:1'h0];
  assign T2904 = T1637[1'h1:1'h1];
  assign T2905 = T1637[2'h2:2'h2];
  assign T2906 = T1637[2'h3:2'h3];
  assign twiddle3_1_80_real = T2909 + T2907;
  assign T2907 = $signed(T2908) / $signed(22'h100000);
  assign T2908 = $signed(31'h383c0315) * $signed(16'h0);
  assign T2909 = {T2912, T2910};
  assign T2910 = $signed(T2911) / $signed(22'h100000);
  assign T2911 = $signed(30'h217193da) * $signed(16'h1);
  assign T2912 = T2910[6'h2d:6'h2d];
  assign T2913 = T1637[3'h4:3'h4];
  assign T2914 = T2773[6'h2e:6'h2e];
  assign T2915 = T1637[3'h6:3'h6];
  assign io_t4_3out_imag = T2916;
  assign T2916 = T2917[4'hf:1'h0];
  assign T2917 = T6853 ? T4895 : T2918;
  assign T2918 = T4894 ? T3871 : T2919;
  assign T2919 = T3870 ? T3458 : T2920;
  assign T2920 = T3457 ? T3215 : T2921;
  assign T2921 = T3214 ? T3074 : T2922;
  assign T2922 = T3073 ? T3001 : T2923;
  assign T2923 = T3000 ? T2964 : T2924;
  assign T2924 = T2963 ? T2945 : T2925;
  assign T2925 = T2942 ? T2933 : twiddle4_3_0_imag;
  assign twiddle4_3_0_imag = T2931 + T2926;
  assign T2926 = {T2929, T2927};
  assign T2927 = $signed(T2928) / $signed(22'h100000);
  assign T2928 = $signed(1'h0) * $signed(16'hffff);
  assign T2929 = T2930 ? 31'h7fffffff : 31'h0;
  assign T2930 = T2927[5'h10:5'h10];
  assign T2931 = $signed(T2932) / $signed(22'h100000);
  assign T2932 = $signed(32'h40000000) * $signed(16'h0);
  assign T2933 = {T2941, twiddle4_3_1_imag};
  assign twiddle4_3_1_imag = T2939 + T2934;
  assign T2934 = {T2937, T2935};
  assign T2935 = $signed(T2936) / $signed(22'h100000);
  assign T2936 = $signed(25'h96cb58) * $signed(16'hffff);
  assign T2937 = T2938 ? 6'h3f : 6'h0;
  assign T2938 = T2935[6'h28:6'h28];
  assign T2939 = $signed(T2940) / $signed(22'h100000);
  assign T2940 = $signed(31'h3fff4e59) * $signed(16'h0);
  assign T2941 = twiddle4_3_1_imag[6'h2e:6'h2e];
  assign T2942 = T2943[1'h0:1'h0];
  assign T2943 = T2944;
  assign T2944 = io_in4[4'h8:1'h0];
  assign T2945 = {T2962, T2946};
  assign T2946 = T2961 ? twiddle4_3_3_imag : twiddle4_3_2_imag;
  assign twiddle4_3_2_imag = T2952 + T2947;
  assign T2947 = {T2950, T2948};
  assign T2948 = $signed(T2949) / $signed(22'h100000);
  assign T2949 = $signed(26'h12d936b) * $signed(16'hffff);
  assign T2950 = T2951 ? 5'h1f : 5'h0;
  assign T2951 = T2948[6'h29:6'h29];
  assign T2952 = $signed(T2953) / $signed(22'h100000);
  assign T2953 = $signed(31'h3ffd3968) * $signed(16'h0);
  assign twiddle4_3_3_imag = T2959 + T2954;
  assign T2954 = {T2957, T2955};
  assign T2955 = $signed(T2956) / $signed(22'h100000);
  assign T2956 = $signed(26'h1c454f4) * $signed(16'hffff);
  assign T2957 = T2958 ? 5'h1f : 5'h0;
  assign T2958 = T2955[6'h29:6'h29];
  assign T2959 = $signed(T2960) / $signed(22'h100000);
  assign T2960 = $signed(31'h3ff9c139) * $signed(16'h0);
  assign T2961 = T2943[1'h0:1'h0];
  assign T2962 = T2946[6'h2e:6'h2e];
  assign T2963 = T2943[1'h1:1'h1];
  assign T2964 = {T2999, T2965};
  assign T2965 = T2998 ? T2982 : T2966;
  assign T2966 = T2981 ? twiddle4_3_5_imag : twiddle4_3_4_imag;
  assign twiddle4_3_4_imag = T2972 + T2967;
  assign T2967 = {T2970, T2968};
  assign T2968 = $signed(T2969) / $signed(22'h100000);
  assign T2969 = $signed(27'h25b0cae) * $signed(16'hffff);
  assign T2970 = T2971 ? 4'hf : 4'h0;
  assign T2971 = T2968[6'h2a:6'h2a];
  assign T2972 = $signed(T2973) / $signed(22'h100000);
  assign T2973 = $signed(31'h3ff4e5df) * $signed(16'h0);
  assign twiddle4_3_5_imag = T2979 + T2974;
  assign T2974 = {T2977, T2975};
  assign T2975 = $signed(T2976) / $signed(22'h100000);
  assign T2976 = $signed(27'h2f1b754) * $signed(16'hffff);
  assign T2977 = T2978 ? 4'hf : 4'h0;
  assign T2978 = T2975[6'h2a:6'h2a];
  assign T2979 = $signed(T2980) / $signed(22'h100000);
  assign T2980 = $signed(31'h3feea776) * $signed(16'h0);
  assign T2981 = T2943[1'h0:1'h0];
  assign T2982 = T2997 ? twiddle4_3_7_imag : twiddle4_3_6_imag;
  assign twiddle4_3_6_imag = T2988 + T2983;
  assign T2983 = {T2986, T2984};
  assign T2984 = $signed(T2985) / $signed(22'h100000);
  assign T2985 = $signed(27'h38851a2) * $signed(16'hffff);
  assign T2986 = T2987 ? 4'hf : 4'h0;
  assign T2987 = T2984[6'h2a:6'h2a];
  assign T2988 = $signed(T2989) / $signed(22'h100000);
  assign T2989 = $signed(31'h3fe7061f) * $signed(16'h0);
  assign twiddle4_3_7_imag = T2995 + T2990;
  assign T2990 = {T2993, T2991};
  assign T2991 = $signed(T2992) / $signed(22'h100000);
  assign T2992 = $signed(28'h41ed853) * $signed(16'hffff);
  assign T2993 = T2994 ? 3'h7 : 3'h0;
  assign T2994 = T2991[6'h2b:6'h2b];
  assign T2995 = $signed(T2996) / $signed(22'h100000);
  assign T2996 = $signed(31'h3fde0205) * $signed(16'h0);
  assign T2997 = T2943[1'h0:1'h0];
  assign T2998 = T2943[1'h1:1'h1];
  assign T2999 = T2965[6'h2e:6'h2e];
  assign T3000 = T2943[2'h2:2'h2];
  assign T3001 = {T3072, T3002};
  assign T3002 = T3071 ? T3037 : T3003;
  assign T3003 = T3036 ? T3020 : T3004;
  assign T3004 = T3019 ? twiddle4_3_9_imag : twiddle4_3_8_imag;
  assign twiddle4_3_8_imag = T3010 + T3005;
  assign T3005 = {T3008, T3006};
  assign T3006 = $signed(T3007) / $signed(22'h100000);
  assign T3007 = $signed(28'h4b54824) * $signed(16'hffff);
  assign T3008 = T3009 ? 3'h7 : 3'h0;
  assign T3009 = T3006[6'h2b:6'h2b];
  assign T3010 = $signed(T3011) / $signed(22'h100000);
  assign T3011 = $signed(31'h3fd39b5a) * $signed(16'h0);
  assign twiddle4_3_9_imag = T3017 + T3012;
  assign T3012 = {T3015, T3013};
  assign T3013 = $signed(T3014) / $signed(22'h100000);
  assign T3014 = $signed(28'h54b9dd2) * $signed(16'hffff);
  assign T3015 = T3016 ? 3'h7 : 3'h0;
  assign T3016 = T3013[6'h2b:6'h2b];
  assign T3017 = $signed(T3018) / $signed(22'h100000);
  assign T3018 = $signed(31'h3fc7d257) * $signed(16'h0);
  assign T3019 = T2943[1'h0:1'h0];
  assign T3020 = T3035 ? twiddle4_3_11_imag : twiddle4_3_10_imag;
  assign twiddle4_3_10_imag = T3026 + T3021;
  assign T3021 = {T3024, T3022};
  assign T3022 = $signed(T3023) / $signed(22'h100000);
  assign T3023 = $signed(28'h5e1d61a) * $signed(16'hffff);
  assign T3024 = T3025 ? 3'h7 : 3'h0;
  assign T3025 = T3022[6'h2b:6'h2b];
  assign T3026 = $signed(T3027) / $signed(22'h100000);
  assign T3027 = $signed(31'h3fbaa73f) * $signed(16'h0);
  assign twiddle4_3_11_imag = T3033 + T3028;
  assign T3028 = {T3031, T3029};
  assign T3029 = $signed(T3030) / $signed(22'h100000);
  assign T3030 = $signed(28'h677edba) * $signed(16'hffff);
  assign T3031 = T3032 ? 3'h7 : 3'h0;
  assign T3032 = T3029[6'h2b:6'h2b];
  assign T3033 = $signed(T3034) / $signed(22'h100000);
  assign T3034 = $signed(31'h3fac1a5b) * $signed(16'h0);
  assign T3035 = T2943[1'h0:1'h0];
  assign T3036 = T2943[1'h1:1'h1];
  assign T3037 = T3070 ? T3054 : T3038;
  assign T3038 = T3053 ? twiddle4_3_13_imag : twiddle4_3_12_imag;
  assign twiddle4_3_12_imag = T3044 + T3039;
  assign T3039 = {T3042, T3040};
  assign T3040 = $signed(T3041) / $signed(22'h100000);
  assign T3041 = $signed(28'h70de171) * $signed(16'hffff);
  assign T3042 = T3043 ? 3'h7 : 3'h0;
  assign T3043 = T3040[6'h2b:6'h2b];
  assign T3044 = $signed(T3045) / $signed(22'h100000);
  assign T3045 = $signed(31'h3f9c2bfa) * $signed(16'h0);
  assign twiddle4_3_13_imag = T3051 + T3046;
  assign T3046 = {T3049, T3047};
  assign T3047 = $signed(T3048) / $signed(22'h100000);
  assign T3048 = $signed(28'h7a3adff) * $signed(16'hffff);
  assign T3049 = T3050 ? 3'h7 : 3'h0;
  assign T3050 = T3047[6'h2b:6'h2b];
  assign T3051 = $signed(T3052) / $signed(22'h100000);
  assign T3052 = $signed(31'h3f8adc76) * $signed(16'h0);
  assign T3053 = T2943[1'h0:1'h0];
  assign T3054 = T3069 ? twiddle4_3_15_imag : twiddle4_3_14_imag;
  assign twiddle4_3_14_imag = T3060 + T3055;
  assign T3055 = {T3058, T3056};
  assign T3056 = $signed(T3057) / $signed(22'h100000);
  assign T3057 = $signed(29'h8395023) * $signed(16'hffff);
  assign T3058 = T3059 ? 2'h3 : 2'h0;
  assign T3059 = T3056[6'h2c:6'h2c];
  assign T3060 = $signed(T3061) / $signed(22'h100000);
  assign T3061 = $signed(31'h3f782c2f) * $signed(16'h0);
  assign twiddle4_3_15_imag = T3067 + T3062;
  assign T3062 = {T3065, T3063};
  assign T3063 = $signed(T3064) / $signed(22'h100000);
  assign T3064 = $signed(29'h8cec4a0) * $signed(16'hffff);
  assign T3065 = T3066 ? 2'h3 : 2'h0;
  assign T3066 = T3063[6'h2c:6'h2c];
  assign T3067 = $signed(T3068) / $signed(22'h100000);
  assign T3068 = $signed(31'h3f641b8d) * $signed(16'h0);
  assign T3069 = T2943[1'h0:1'h0];
  assign T3070 = T2943[1'h1:1'h1];
  assign T3071 = T2943[2'h2:2'h2];
  assign T3072 = T3002[6'h2e:6'h2e];
  assign T3073 = T2943[2'h3:2'h3];
  assign T3074 = {T3213, T3075};
  assign T3075 = T3212 ? T3146 : T3076;
  assign T3076 = T3145 ? T3111 : T3077;
  assign T3077 = T3110 ? T3094 : T3078;
  assign T3078 = T3093 ? twiddle4_3_17_imag : twiddle4_3_16_imag;
  assign twiddle4_3_16_imag = T3084 + T3079;
  assign T3079 = {T3082, T3080};
  assign T3080 = $signed(T3081) / $signed(22'h100000);
  assign T3081 = $signed(29'h9640837) * $signed(16'hffff);
  assign T3082 = T3083 ? 2'h3 : 2'h0;
  assign T3083 = T3080[6'h2c:6'h2c];
  assign T3084 = $signed(T3085) / $signed(22'h100000);
  assign T3085 = $signed(31'h3f4eaafe) * $signed(16'h0);
  assign twiddle4_3_17_imag = T3091 + T3086;
  assign T3086 = {T3089, T3087};
  assign T3087 = $signed(T3088) / $signed(22'h100000);
  assign T3088 = $signed(29'h9f917ab) * $signed(16'hffff);
  assign T3089 = T3090 ? 2'h3 : 2'h0;
  assign T3090 = T3087[6'h2c:6'h2c];
  assign T3091 = $signed(T3092) / $signed(22'h100000);
  assign T3092 = $signed(31'h3f37daf9) * $signed(16'h0);
  assign T3093 = T2943[1'h0:1'h0];
  assign T3094 = T3109 ? twiddle4_3_19_imag : twiddle4_3_18_imag;
  assign twiddle4_3_18_imag = T3100 + T3095;
  assign T3095 = {T3098, T3096};
  assign T3096 = $signed(T3097) / $signed(22'h100000);
  assign T3097 = $signed(29'ha8defc2) * $signed(16'hffff);
  assign T3098 = T3099 ? 2'h3 : 2'h0;
  assign T3099 = T3096[6'h2c:6'h2c];
  assign T3100 = $signed(T3101) / $signed(22'h100000);
  assign T3101 = $signed(31'h3f1fabff) * $signed(16'h0);
  assign twiddle4_3_19_imag = T3107 + T3102;
  assign T3102 = {T3105, T3103};
  assign T3103 = $signed(T3104) / $signed(22'h100000);
  assign T3104 = $signed(29'hb228d41) * $signed(16'hffff);
  assign T3105 = T3106 ? 2'h3 : 2'h0;
  assign T3106 = T3103[6'h2c:6'h2c];
  assign T3107 = $signed(T3108) / $signed(22'h100000);
  assign T3108 = $signed(31'h3f061e94) * $signed(16'h0);
  assign T3109 = T2943[1'h0:1'h0];
  assign T3110 = T2943[1'h1:1'h1];
  assign T3111 = T3144 ? T3128 : T3112;
  assign T3112 = T3127 ? twiddle4_3_21_imag : twiddle4_3_20_imag;
  assign twiddle4_3_20_imag = T3118 + T3113;
  assign T3113 = {T3116, T3114};
  assign T3114 = $signed(T3115) / $signed(22'h100000);
  assign T3115 = $signed(29'hbb6ecef) * $signed(16'hffff);
  assign T3116 = T3117 ? 2'h3 : 2'h0;
  assign T3117 = T3114[6'h2c:6'h2c];
  assign T3118 = $signed(T3119) / $signed(22'h100000);
  assign T3119 = $signed(31'h3eeb3347) * $signed(16'h0);
  assign twiddle4_3_21_imag = T3125 + T3120;
  assign T3120 = {T3123, T3121};
  assign T3121 = $signed(T3122) / $signed(22'h100000);
  assign T3122 = $signed(29'hc4b0b93) * $signed(16'hffff);
  assign T3123 = T3124 ? 2'h3 : 2'h0;
  assign T3124 = T3121[6'h2c:6'h2c];
  assign T3125 = $signed(T3126) / $signed(22'h100000);
  assign T3126 = $signed(31'h3eceeaad) * $signed(16'h0);
  assign T3127 = T2943[1'h0:1'h0];
  assign T3128 = T3143 ? twiddle4_3_23_imag : twiddle4_3_22_imag;
  assign twiddle4_3_22_imag = T3134 + T3129;
  assign T3129 = {T3132, T3130};
  assign T3130 = $signed(T3131) / $signed(22'h100000);
  assign T3131 = $signed(29'hcdee5f9) * $signed(16'hffff);
  assign T3132 = T3133 ? 2'h3 : 2'h0;
  assign T3133 = T3130[6'h2c:6'h2c];
  assign T3134 = $signed(T3135) / $signed(22'h100000);
  assign T3135 = $signed(31'h3eb14562) * $signed(16'h0);
  assign twiddle4_3_23_imag = T3141 + T3136;
  assign T3136 = {T3139, T3137};
  assign T3137 = $signed(T3138) / $signed(22'h100000);
  assign T3138 = $signed(29'hd7278ea) * $signed(16'hffff);
  assign T3139 = T3140 ? 2'h3 : 2'h0;
  assign T3140 = T3137[6'h2c:6'h2c];
  assign T3141 = $signed(T3142) / $signed(22'h100000);
  assign T3142 = $signed(31'h3e92440d) * $signed(16'h0);
  assign T3143 = T2943[1'h0:1'h0];
  assign T3144 = T2943[1'h1:1'h1];
  assign T3145 = T2943[2'h2:2'h2];
  assign T3146 = T3211 ? T3181 : T3147;
  assign T3147 = T3180 ? T3164 : T3148;
  assign T3148 = T3163 ? twiddle4_3_25_imag : twiddle4_3_24_imag;
  assign twiddle4_3_24_imag = T3154 + T3149;
  assign T3149 = {T3152, T3150};
  assign T3150 = $signed(T3151) / $signed(22'h100000);
  assign T3151 = $signed(29'he05c135) * $signed(16'hffff);
  assign T3152 = T3153 ? 2'h3 : 2'h0;
  assign T3153 = T3150[6'h2c:6'h2c];
  assign T3154 = $signed(T3155) / $signed(22'h100000);
  assign T3155 = $signed(31'h3e71e758) * $signed(16'h0);
  assign twiddle4_3_25_imag = T3161 + T3156;
  assign T3156 = {T3159, T3157};
  assign T3157 = $signed(T3158) / $signed(22'h100000);
  assign T3158 = $signed(29'he98bba6) * $signed(16'hffff);
  assign T3159 = T3160 ? 2'h3 : 2'h0;
  assign T3160 = T3157[6'h2c:6'h2c];
  assign T3161 = $signed(T3162) / $signed(22'h100000);
  assign T3162 = $signed(31'h3e502ff8) * $signed(16'h0);
  assign T3163 = T2943[1'h0:1'h0];
  assign T3164 = T3179 ? twiddle4_3_27_imag : twiddle4_3_26_imag;
  assign twiddle4_3_26_imag = T3170 + T3165;
  assign T3165 = {T3168, T3166};
  assign T3166 = $signed(T3167) / $signed(22'h100000);
  assign T3167 = $signed(29'hf2b650f) * $signed(16'hffff);
  assign T3168 = T3169 ? 2'h3 : 2'h0;
  assign T3169 = T3166[6'h2c:6'h2c];
  assign T3170 = $signed(T3171) / $signed(22'h100000);
  assign T3171 = $signed(31'h3e2d1ea7) * $signed(16'h0);
  assign twiddle4_3_27_imag = T3177 + T3172;
  assign T3172 = {T3175, T3173};
  assign T3173 = $signed(T3174) / $signed(22'h100000);
  assign T3174 = $signed(29'hfbdba40) * $signed(16'hffff);
  assign T3175 = T3176 ? 2'h3 : 2'h0;
  assign T3176 = T3173[6'h2c:6'h2c];
  assign T3177 = $signed(T3178) / $signed(22'h100000);
  assign T3178 = $signed(31'h3e08b429) * $signed(16'h0);
  assign T3179 = T2943[1'h0:1'h0];
  assign T3180 = T2943[1'h1:1'h1];
  assign T3181 = T3210 ? T3196 : T3182;
  assign T3182 = T3195 ? twiddle4_3_29_imag : twiddle4_3_28_imag;
  assign twiddle4_3_28_imag = T3187 + T3183;
  assign T3183 = {T3186, T3184};
  assign T3184 = $signed(T3185) / $signed(22'h100000);
  assign T3185 = $signed(30'h104fb80e) * $signed(16'hffff);
  assign T3186 = T3184[6'h2d:6'h2d];
  assign T3187 = $signed(T3188) / $signed(22'h100000);
  assign T3188 = $signed(31'h3de2f147) * $signed(16'h0);
  assign twiddle4_3_29_imag = T3193 + T3189;
  assign T3189 = {T3192, T3190};
  assign T3190 = $signed(T3191) / $signed(22'h100000);
  assign T3191 = $signed(30'h10e15b4e) * $signed(16'hffff);
  assign T3192 = T3190[6'h2d:6'h2d];
  assign T3193 = $signed(T3194) / $signed(22'h100000);
  assign T3194 = $signed(31'h3dbbd6d4) * $signed(16'h0);
  assign T3195 = T2943[1'h0:1'h0];
  assign T3196 = T3209 ? twiddle4_3_31_imag : twiddle4_3_30_imag;
  assign twiddle4_3_30_imag = T3201 + T3197;
  assign T3197 = {T3200, T3198};
  assign T3198 = $signed(T3199) / $signed(22'h100000);
  assign T3199 = $signed(30'h1172a0d7) * $signed(16'hffff);
  assign T3200 = T3198[6'h2d:6'h2d];
  assign T3201 = $signed(T3202) / $signed(22'h100000);
  assign T3202 = $signed(31'h3d9365a7) * $signed(16'h0);
  assign twiddle4_3_31_imag = T3207 + T3203;
  assign T3203 = {T3206, T3204};
  assign T3204 = $signed(T3205) / $signed(22'h100000);
  assign T3205 = $signed(30'h12038583) * $signed(16'hffff);
  assign T3206 = T3204[6'h2d:6'h2d];
  assign T3207 = $signed(T3208) / $signed(22'h100000);
  assign T3208 = $signed(31'h3d699ea2) * $signed(16'h0);
  assign T3209 = T2943[1'h0:1'h0];
  assign T3210 = T2943[1'h1:1'h1];
  assign T3211 = T2943[2'h2:2'h2];
  assign T3212 = T2943[2'h3:2'h3];
  assign T3213 = T3075[6'h2e:6'h2e];
  assign T3214 = T2943[3'h4:3'h4];
  assign T3215 = {T3456, T3216};
  assign T3216 = T3455 ? T3343 : T3217;
  assign T3217 = T3342 ? T3280 : T3218;
  assign T3218 = T3279 ? T3249 : T3219;
  assign T3219 = T3248 ? T3234 : T3220;
  assign T3220 = T3233 ? twiddle4_3_33_imag : twiddle4_3_32_imag;
  assign twiddle4_3_32_imag = T3225 + T3221;
  assign T3221 = {T3224, T3222};
  assign T3222 = $signed(T3223) / $signed(22'h100000);
  assign T3223 = $signed(30'h1294062e) * $signed(16'hffff);
  assign T3224 = T3222[6'h2d:6'h2d];
  assign T3225 = $signed(T3226) / $signed(22'h100000);
  assign T3226 = $signed(31'h3d3e82ad) * $signed(16'h0);
  assign twiddle4_3_33_imag = T3231 + T3227;
  assign T3227 = {T3230, T3228};
  assign T3228 = $signed(T3229) / $signed(22'h100000);
  assign T3229 = $signed(30'h13241fb6) * $signed(16'hffff);
  assign T3230 = T3228[6'h2d:6'h2d];
  assign T3231 = $signed(T3232) / $signed(22'h100000);
  assign T3232 = $signed(31'h3d1212b7) * $signed(16'h0);
  assign T3233 = T2943[1'h0:1'h0];
  assign T3234 = T3247 ? twiddle4_3_35_imag : twiddle4_3_34_imag;
  assign twiddle4_3_34_imag = T3239 + T3235;
  assign T3235 = {T3238, T3236};
  assign T3236 = $signed(T3237) / $signed(22'h100000);
  assign T3237 = $signed(30'h13b3cefa) * $signed(16'hffff);
  assign T3238 = T3236[6'h2d:6'h2d];
  assign T3239 = $signed(T3240) / $signed(22'h100000);
  assign T3240 = $signed(31'h3ce44fb6) * $signed(16'h0);
  assign twiddle4_3_35_imag = T3245 + T3241;
  assign T3241 = {T3244, T3242};
  assign T3242 = $signed(T3243) / $signed(22'h100000);
  assign T3243 = $signed(30'h144310dc) * $signed(16'hffff);
  assign T3244 = T3242[6'h2d:6'h2d];
  assign T3245 = $signed(T3246) / $signed(22'h100000);
  assign T3246 = $signed(31'h3cb53aaa) * $signed(16'h0);
  assign T3247 = T2943[1'h0:1'h0];
  assign T3248 = T2943[1'h1:1'h1];
  assign T3249 = T3278 ? T3264 : T3250;
  assign T3250 = T3263 ? twiddle4_3_37_imag : twiddle4_3_36_imag;
  assign twiddle4_3_36_imag = T3255 + T3251;
  assign T3251 = {T3254, T3252};
  assign T3252 = $signed(T3253) / $signed(22'h100000);
  assign T3253 = $signed(30'h14d1e242) * $signed(16'hffff);
  assign T3254 = T3252[6'h2d:6'h2d];
  assign T3255 = $signed(T3256) / $signed(22'h100000);
  assign T3256 = $signed(31'h3c84d496) * $signed(16'h0);
  assign twiddle4_3_37_imag = T3261 + T3257;
  assign T3257 = {T3260, T3258};
  assign T3258 = $signed(T3259) / $signed(22'h100000);
  assign T3259 = $signed(30'h15604012) * $signed(16'hffff);
  assign T3260 = T3258[6'h2d:6'h2d];
  assign T3261 = $signed(T3262) / $signed(22'h100000);
  assign T3262 = $signed(31'h3c531e88) * $signed(16'h0);
  assign T3263 = T2943[1'h0:1'h0];
  assign T3264 = T3277 ? twiddle4_3_39_imag : twiddle4_3_38_imag;
  assign twiddle4_3_38_imag = T3269 + T3265;
  assign T3265 = {T3268, T3266};
  assign T3266 = $signed(T3267) / $signed(22'h100000);
  assign T3267 = $signed(30'h15ee2737) * $signed(16'hffff);
  assign T3268 = T3266[6'h2d:6'h2d];
  assign T3269 = $signed(T3270) / $signed(22'h100000);
  assign T3270 = $signed(31'h3c201994) * $signed(16'h0);
  assign twiddle4_3_39_imag = T3275 + T3271;
  assign T3271 = {T3274, T3272};
  assign T3272 = $signed(T3273) / $signed(22'h100000);
  assign T3273 = $signed(30'h167b949c) * $signed(16'hffff);
  assign T3274 = T3272[6'h2d:6'h2d];
  assign T3275 = $signed(T3276) / $signed(22'h100000);
  assign T3276 = $signed(31'h3bebc6d5) * $signed(16'h0);
  assign T3277 = T2943[1'h0:1'h0];
  assign T3278 = T2943[1'h1:1'h1];
  assign T3279 = T2943[2'h2:2'h2];
  assign T3280 = T3341 ? T3311 : T3281;
  assign T3281 = T3310 ? T3296 : T3282;
  assign T3282 = T3295 ? twiddle4_3_41_imag : twiddle4_3_40_imag;
  assign twiddle4_3_40_imag = T3287 + T3283;
  assign T3283 = {T3286, T3284};
  assign T3284 = $signed(T3285) / $signed(22'h100000);
  assign T3285 = $signed(30'h17088530) * $signed(16'hffff);
  assign T3286 = T3284[6'h2d:6'h2d];
  assign T3287 = $signed(T3288) / $signed(22'h100000);
  assign T3288 = $signed(31'h3bb6276d) * $signed(16'h0);
  assign twiddle4_3_41_imag = T3293 + T3289;
  assign T3289 = {T3292, T3290};
  assign T3290 = $signed(T3291) / $signed(22'h100000);
  assign T3291 = $signed(30'h1794f5e6) * $signed(16'hffff);
  assign T3292 = T3290[6'h2d:6'h2d];
  assign T3293 = $signed(T3294) / $signed(22'h100000);
  assign T3294 = $signed(31'h3b7f3c87) * $signed(16'h0);
  assign T3295 = T2943[1'h0:1'h0];
  assign T3296 = T3309 ? twiddle4_3_43_imag : twiddle4_3_42_imag;
  assign twiddle4_3_42_imag = T3301 + T3297;
  assign T3297 = {T3300, T3298};
  assign T3298 = $signed(T3299) / $signed(22'h100000);
  assign T3299 = $signed(30'h1820e3b0) * $signed(16'hffff);
  assign T3300 = T3298[6'h2d:6'h2d];
  assign T3301 = $signed(T3302) / $signed(22'h100000);
  assign T3302 = $signed(31'h3b470752) * $signed(16'h0);
  assign twiddle4_3_43_imag = T3307 + T3303;
  assign T3303 = {T3306, T3304};
  assign T3304 = $signed(T3305) / $signed(22'h100000);
  assign T3305 = $signed(30'h18ac4b86) * $signed(16'hffff);
  assign T3306 = T3304[6'h2d:6'h2d];
  assign T3307 = $signed(T3308) / $signed(22'h100000);
  assign T3308 = $signed(31'h3b0d8908) * $signed(16'h0);
  assign T3309 = T2943[1'h0:1'h0];
  assign T3310 = T2943[1'h1:1'h1];
  assign T3311 = T3340 ? T3326 : T3312;
  assign T3312 = T3325 ? twiddle4_3_45_imag : twiddle4_3_44_imag;
  assign twiddle4_3_44_imag = T3317 + T3313;
  assign T3313 = {T3316, T3314};
  assign T3314 = $signed(T3315) / $signed(22'h100000);
  assign T3315 = $signed(30'h19372a63) * $signed(16'hffff);
  assign T3316 = T3314[6'h2d:6'h2d];
  assign T3317 = $signed(T3318) / $signed(22'h100000);
  assign T3318 = $signed(31'h3ad2c2e7) * $signed(16'h0);
  assign twiddle4_3_45_imag = T3323 + T3319;
  assign T3319 = {T3322, T3320};
  assign T3320 = $signed(T3321) / $signed(22'h100000);
  assign T3321 = $signed(30'h19c17d44) * $signed(16'hffff);
  assign T3322 = T3320[6'h2d:6'h2d];
  assign T3323 = $signed(T3324) / $signed(22'h100000);
  assign T3324 = $signed(31'h3a96b636) * $signed(16'h0);
  assign T3325 = T2943[1'h0:1'h0];
  assign T3326 = T3339 ? twiddle4_3_47_imag : twiddle4_3_46_imag;
  assign twiddle4_3_46_imag = T3331 + T3327;
  assign T3327 = {T3330, T3328};
  assign T3328 = $signed(T3329) / $signed(22'h100000);
  assign T3329 = $signed(30'h1a4b4127) * $signed(16'hffff);
  assign T3330 = T3328[6'h2d:6'h2d];
  assign T3331 = $signed(T3332) / $signed(22'h100000);
  assign T3332 = $signed(31'h3a596441) * $signed(16'h0);
  assign twiddle4_3_47_imag = T3337 + T3333;
  assign T3333 = {T3336, T3334};
  assign T3334 = $signed(T3335) / $signed(22'h100000);
  assign T3335 = $signed(30'h1ad47312) * $signed(16'hffff);
  assign T3336 = T3334[6'h2d:6'h2d];
  assign T3337 = $signed(T3338) / $signed(22'h100000);
  assign T3338 = $signed(31'h3a1ace5e) * $signed(16'h0);
  assign T3339 = T2943[1'h0:1'h0];
  assign T3340 = T2943[1'h1:1'h1];
  assign T3341 = T2943[2'h2:2'h2];
  assign T3342 = T2943[2'h3:2'h3];
  assign T3343 = T3454 ? T3406 : T3344;
  assign T3344 = T3405 ? T3375 : T3345;
  assign T3345 = T3374 ? T3360 : T3346;
  assign T3346 = T3359 ? twiddle4_3_49_imag : twiddle4_3_48_imag;
  assign twiddle4_3_48_imag = T3351 + T3347;
  assign T3347 = {T3350, T3348};
  assign T3348 = $signed(T3349) / $signed(22'h100000);
  assign T3349 = $signed(30'h1b5d1009) * $signed(16'hffff);
  assign T3350 = T3348[6'h2d:6'h2d];
  assign T3351 = $signed(T3352) / $signed(22'h100000);
  assign T3352 = $signed(31'h39daf5e8) * $signed(16'h0);
  assign twiddle4_3_49_imag = T3357 + T3353;
  assign T3353 = {T3356, T3354};
  assign T3354 = $signed(T3355) / $signed(22'h100000);
  assign T3355 = $signed(30'h1be51517) * $signed(16'hffff);
  assign T3356 = T3354[6'h2d:6'h2d];
  assign T3357 = $signed(T3358) / $signed(22'h100000);
  assign T3358 = $signed(31'h3999dc41) * $signed(16'h0);
  assign T3359 = T2943[1'h0:1'h0];
  assign T3360 = T3373 ? twiddle4_3_51_imag : twiddle4_3_50_imag;
  assign twiddle4_3_50_imag = T3365 + T3361;
  assign T3361 = {T3364, T3362};
  assign T3362 = $signed(T3363) / $signed(22'h100000);
  assign T3363 = $signed(30'h1c6c7f49) * $signed(16'hffff);
  assign T3364 = T3362[6'h2d:6'h2d];
  assign T3365 = $signed(T3366) / $signed(22'h100000);
  assign T3366 = $signed(31'h395782d3) * $signed(16'h0);
  assign twiddle4_3_51_imag = T3371 + T3367;
  assign T3367 = {T3370, T3368};
  assign T3368 = $signed(T3369) / $signed(22'h100000);
  assign T3369 = $signed(30'h1cf34bae) * $signed(16'hffff);
  assign T3370 = T3368[6'h2d:6'h2d];
  assign T3371 = $signed(T3372) / $signed(22'h100000);
  assign T3372 = $signed(31'h3913eb0e) * $signed(16'h0);
  assign T3373 = T2943[1'h0:1'h0];
  assign T3374 = T2943[1'h1:1'h1];
  assign T3375 = T3404 ? T3390 : T3376;
  assign T3376 = T3389 ? twiddle4_3_53_imag : twiddle4_3_52_imag;
  assign twiddle4_3_52_imag = T3381 + T3377;
  assign T3377 = {T3380, T3378};
  assign T3378 = $signed(T3379) / $signed(22'h100000);
  assign T3379 = $signed(30'h1d79775b) * $signed(16'hffff);
  assign T3380 = T3378[6'h2d:6'h2d];
  assign T3381 = $signed(T3382) / $signed(22'h100000);
  assign T3382 = $signed(31'h38cf1669) * $signed(16'h0);
  assign twiddle4_3_53_imag = T3387 + T3383;
  assign T3383 = {T3386, T3384};
  assign T3384 = $signed(T3385) / $signed(22'h100000);
  assign T3385 = $signed(30'h1dfeff66) * $signed(16'hffff);
  assign T3386 = T3384[6'h2d:6'h2d];
  assign T3387 = $signed(T3388) / $signed(22'h100000);
  assign T3388 = $signed(31'h38890662) * $signed(16'h0);
  assign T3389 = T2943[1'h0:1'h0];
  assign T3390 = T3403 ? twiddle4_3_55_imag : twiddle4_3_54_imag;
  assign twiddle4_3_54_imag = T3395 + T3391;
  assign T3391 = {T3394, T3392};
  assign T3392 = $signed(T3393) / $signed(22'h100000);
  assign T3393 = $signed(30'h1e83e0ea) * $signed(16'hffff);
  assign T3394 = T3392[6'h2d:6'h2d];
  assign T3395 = $signed(T3396) / $signed(22'h100000);
  assign T3396 = $signed(31'h3841bc7f) * $signed(16'h0);
  assign twiddle4_3_55_imag = T3401 + T3397;
  assign T3397 = {T3400, T3398};
  assign T3398 = $signed(T3399) / $signed(22'h100000);
  assign T3399 = $signed(30'h1f081906) * $signed(16'hffff);
  assign T3400 = T3398[6'h2d:6'h2d];
  assign T3401 = $signed(T3402) / $signed(22'h100000);
  assign T3402 = $signed(31'h37f93a4b) * $signed(16'h0);
  assign T3403 = T2943[1'h0:1'h0];
  assign T3404 = T2943[1'h1:1'h1];
  assign T3405 = T2943[2'h2:2'h2];
  assign T3406 = T3453 ? T3431 : T3407;
  assign T3407 = T3430 ? T3420 : T3408;
  assign T3408 = T3419 ? twiddle4_3_57_imag : twiddle4_3_56_imag;
  assign twiddle4_3_56_imag = T3413 + T3409;
  assign T3409 = {T3412, T3410};
  assign T3410 = $signed(T3411) / $signed(22'h100000);
  assign T3411 = $signed(30'h1f8ba4db) * $signed(16'hffff);
  assign T3412 = T3410[6'h2d:6'h2d];
  assign T3413 = $signed(T3414) / $signed(22'h100000);
  assign T3414 = $signed(31'h37af8158) * $signed(16'h0);
  assign twiddle4_3_57_imag = T3417 + T3415;
  assign T3415 = $signed(T3416) / $signed(22'h100000);
  assign T3416 = $signed(31'h200e8190) * $signed(16'hffff);
  assign T3417 = $signed(T3418) / $signed(22'h100000);
  assign T3418 = $signed(31'h37649341) * $signed(16'h0);
  assign T3419 = T2943[1'h0:1'h0];
  assign T3420 = T3429 ? twiddle4_3_59_imag : twiddle4_3_58_imag;
  assign twiddle4_3_58_imag = T3423 + T3421;
  assign T3421 = $signed(T3422) / $signed(22'h100000);
  assign T3422 = $signed(31'h2090ac4d) * $signed(16'hffff);
  assign T3423 = $signed(T3424) / $signed(22'h100000);
  assign T3424 = $signed(31'h371871a4) * $signed(16'h0);
  assign twiddle4_3_59_imag = T3427 + T3425;
  assign T3425 = $signed(T3426) / $signed(22'h100000);
  assign T3426 = $signed(31'h21122240) * $signed(16'hffff);
  assign T3427 = $signed(T3428) / $signed(22'h100000);
  assign T3428 = $signed(31'h36cb1e29) * $signed(16'h0);
  assign T3429 = T2943[1'h0:1'h0];
  assign T3430 = T2943[1'h1:1'h1];
  assign T3431 = T3452 ? T3442 : T3432;
  assign T3432 = T3441 ? twiddle4_3_61_imag : twiddle4_3_60_imag;
  assign twiddle4_3_60_imag = T3435 + T3433;
  assign T3433 = $signed(T3434) / $signed(22'h100000);
  assign T3434 = $signed(31'h2192e09a) * $signed(16'hffff);
  assign T3435 = $signed(T3436) / $signed(22'h100000);
  assign T3436 = $signed(31'h367c9a7d) * $signed(16'h0);
  assign twiddle4_3_61_imag = T3439 + T3437;
  assign T3437 = $signed(T3438) / $signed(22'h100000);
  assign T3438 = $signed(31'h2212e491) * $signed(16'hffff);
  assign T3439 = $signed(T3440) / $signed(22'h100000);
  assign T3440 = $signed(31'h362ce854) * $signed(16'h0);
  assign T3441 = T2943[1'h0:1'h0];
  assign T3442 = T3451 ? twiddle4_3_63_imag : twiddle4_3_62_imag;
  assign twiddle4_3_62_imag = T3445 + T3443;
  assign T3443 = $signed(T3444) / $signed(22'h100000);
  assign T3444 = $signed(31'h22922b5e) * $signed(16'hffff);
  assign T3445 = $signed(T3446) / $signed(22'h100000);
  assign T3446 = $signed(31'h35dc0968) * $signed(16'h0);
  assign twiddle4_3_63_imag = T3449 + T3447;
  assign T3447 = $signed(T3448) / $signed(22'h100000);
  assign T3448 = $signed(31'h2310b23e) * $signed(16'hffff);
  assign T3449 = $signed(T3450) / $signed(22'h100000);
  assign T3450 = $signed(31'h3589ff7a) * $signed(16'h0);
  assign T3451 = T2943[1'h0:1'h0];
  assign T3452 = T2943[1'h1:1'h1];
  assign T3453 = T2943[2'h2:2'h2];
  assign T3454 = T2943[2'h3:2'h3];
  assign T3455 = T2943[3'h4:3'h4];
  assign T3456 = T3216[6'h2e:6'h2e];
  assign T3457 = T2943[3'h5:3'h5];
  assign T3458 = {T3869, T3459};
  assign T3459 = T3868 ? T3650 : T3460;
  assign T3460 = T3649 ? T3555 : T3461;
  assign T3461 = T3554 ? T3508 : T3462;
  assign T3462 = T3507 ? T3485 : T3463;
  assign T3463 = T3484 ? T3474 : T3464;
  assign T3464 = T3473 ? twiddle4_3_65_imag : twiddle4_3_64_imag;
  assign twiddle4_3_64_imag = T3467 + T3465;
  assign T3465 = $signed(T3466) / $signed(22'h100000);
  assign T3466 = $signed(31'h238e7673) * $signed(16'hffff);
  assign T3467 = $signed(T3468) / $signed(22'h100000);
  assign T3468 = $signed(31'h3536cc52) * $signed(16'h0);
  assign twiddle4_3_65_imag = T3471 + T3469;
  assign T3469 = $signed(T3470) / $signed(22'h100000);
  assign T3470 = $signed(31'h240b7542) * $signed(16'hffff);
  assign T3471 = $signed(T3472) / $signed(22'h100000);
  assign T3472 = $signed(31'h34e271bd) * $signed(16'h0);
  assign T3473 = T2943[1'h0:1'h0];
  assign T3474 = T3483 ? twiddle4_3_67_imag : twiddle4_3_66_imag;
  assign twiddle4_3_66_imag = T3477 + T3475;
  assign T3475 = $signed(T3476) / $signed(22'h100000);
  assign T3476 = $signed(31'h2487abf7) * $signed(16'hffff);
  assign T3477 = $signed(T3478) / $signed(22'h100000);
  assign T3478 = $signed(31'h348cf190) * $signed(16'h0);
  assign twiddle4_3_67_imag = T3481 + T3479;
  assign T3479 = $signed(T3480) / $signed(22'h100000);
  assign T3480 = $signed(31'h250317de) * $signed(16'hffff);
  assign T3481 = $signed(T3482) / $signed(22'h100000);
  assign T3482 = $signed(31'h34364da5) * $signed(16'h0);
  assign T3483 = T2943[1'h0:1'h0];
  assign T3484 = T2943[1'h1:1'h1];
  assign T3485 = T3506 ? T3496 : T3486;
  assign T3486 = T3495 ? twiddle4_3_69_imag : twiddle4_3_68_imag;
  assign twiddle4_3_68_imag = T3489 + T3487;
  assign T3487 = $signed(T3488) / $signed(22'h100000);
  assign T3488 = $signed(31'h257db64b) * $signed(16'hffff);
  assign T3489 = $signed(T3490) / $signed(22'h100000);
  assign T3490 = $signed(31'h33de87de) * $signed(16'h0);
  assign twiddle4_3_69_imag = T3493 + T3491;
  assign T3491 = $signed(T3492) / $signed(22'h100000);
  assign T3492 = $signed(31'h25f78496) * $signed(16'hffff);
  assign T3493 = $signed(T3494) / $signed(22'h100000);
  assign T3494 = $signed(31'h3385a221) * $signed(16'h0);
  assign T3495 = T2943[1'h0:1'h0];
  assign T3496 = T3505 ? twiddle4_3_71_imag : twiddle4_3_70_imag;
  assign twiddle4_3_70_imag = T3499 + T3497;
  assign T3497 = $signed(T3498) / $signed(22'h100000);
  assign T3498 = $signed(31'h2670801a) * $signed(16'hffff);
  assign T3499 = $signed(T3500) / $signed(22'h100000);
  assign T3500 = $signed(31'h332b9e5d) * $signed(16'h0);
  assign twiddle4_3_71_imag = T3503 + T3501;
  assign T3501 = $signed(T3502) / $signed(22'h100000);
  assign T3502 = $signed(31'h26e8a637) * $signed(16'hffff);
  assign T3503 = $signed(T3504) / $signed(22'h100000);
  assign T3504 = $signed(31'h32d07e85) * $signed(16'h0);
  assign T3505 = T2943[1'h0:1'h0];
  assign T3506 = T2943[1'h1:1'h1];
  assign T3507 = T2943[2'h2:2'h2];
  assign T3508 = T3553 ? T3531 : T3509;
  assign T3509 = T3530 ? T3520 : T3510;
  assign T3510 = T3519 ? twiddle4_3_73_imag : twiddle4_3_72_imag;
  assign twiddle4_3_72_imag = T3513 + T3511;
  assign T3511 = $signed(T3512) / $signed(22'h100000);
  assign T3512 = $signed(31'h275ff452) * $signed(16'hffff);
  assign T3513 = $signed(T3514) / $signed(22'h100000);
  assign T3514 = $signed(31'h32744493) * $signed(16'h0);
  assign twiddle4_3_73_imag = T3517 + T3515;
  assign T3515 = $signed(T3516) / $signed(22'h100000);
  assign T3516 = $signed(31'h27d667d5) * $signed(16'hffff);
  assign T3517 = $signed(T3518) / $signed(22'h100000);
  assign T3518 = $signed(31'h3216f286) * $signed(16'h0);
  assign T3519 = T2943[1'h0:1'h0];
  assign T3520 = T3529 ? twiddle4_3_75_imag : twiddle4_3_74_imag;
  assign twiddle4_3_74_imag = T3523 + T3521;
  assign T3521 = $signed(T3522) / $signed(22'h100000);
  assign T3522 = $signed(31'h284bfe2f) * $signed(16'hffff);
  assign T3523 = $signed(T3524) / $signed(22'h100000);
  assign T3524 = $signed(31'h31b88a66) * $signed(16'h0);
  assign twiddle4_3_75_imag = T3527 + T3525;
  assign T3525 = $signed(T3526) / $signed(22'h100000);
  assign T3526 = $signed(31'h28c0b4d2) * $signed(16'hffff);
  assign T3527 = $signed(T3528) / $signed(22'h100000);
  assign T3528 = $signed(31'h31590e3d) * $signed(16'h0);
  assign T3529 = T2943[1'h0:1'h0];
  assign T3530 = T2943[1'h1:1'h1];
  assign T3531 = T3552 ? T3542 : T3532;
  assign T3532 = T3541 ? twiddle4_3_77_imag : twiddle4_3_76_imag;
  assign twiddle4_3_76_imag = T3535 + T3533;
  assign T3533 = $signed(T3534) / $signed(22'h100000);
  assign T3534 = $signed(31'h29348937) * $signed(16'hffff);
  assign T3535 = $signed(T3536) / $signed(22'h100000);
  assign T3536 = $signed(31'h30f8801f) * $signed(16'h0);
  assign twiddle4_3_77_imag = T3539 + T3537;
  assign T3537 = $signed(T3538) / $signed(22'h100000);
  assign T3538 = $signed(31'h29a778da) * $signed(16'hffff);
  assign T3539 = $signed(T3540) / $signed(22'h100000);
  assign T3540 = $signed(31'h3096e223) * $signed(16'h0);
  assign T3541 = T2943[1'h0:1'h0];
  assign T3542 = T3551 ? twiddle4_3_79_imag : twiddle4_3_78_imag;
  assign twiddle4_3_78_imag = T3545 + T3543;
  assign T3543 = $signed(T3544) / $signed(22'h100000);
  assign T3544 = $signed(31'h2a19813e) * $signed(16'hffff);
  assign T3545 = $signed(T3546) / $signed(22'h100000);
  assign T3546 = $signed(31'h30343667) * $signed(16'h0);
  assign twiddle4_3_79_imag = T3549 + T3547;
  assign T3547 = $signed(T3548) / $signed(22'h100000);
  assign T3548 = $signed(31'h2a8a9fea) * $signed(16'hffff);
  assign T3549 = $signed(T3550) / $signed(22'h100000);
  assign T3550 = $signed(31'h2fd07f0f) * $signed(16'h0);
  assign T3551 = T2943[1'h0:1'h0];
  assign T3552 = T2943[1'h1:1'h1];
  assign T3553 = T2943[2'h2:2'h2];
  assign T3554 = T2943[2'h3:2'h3];
  assign T3555 = T3648 ? T3602 : T3556;
  assign T3556 = T3601 ? T3579 : T3557;
  assign T3557 = T3578 ? T3568 : T3558;
  assign T3558 = T3567 ? twiddle4_3_81_imag : twiddle4_3_80_imag;
  assign twiddle4_3_80_imag = T3561 + T3559;
  assign T3559 = $signed(T3560) / $signed(22'h100000);
  assign T3560 = $signed(31'h2afad269) * $signed(16'hffff);
  assign T3561 = $signed(T3562) / $signed(22'h100000);
  assign T3562 = $signed(31'h2f6bbe44) * $signed(16'h0);
  assign twiddle4_3_81_imag = T3565 + T3563;
  assign T3563 = $signed(T3564) / $signed(22'h100000);
  assign T3564 = $signed(31'h2b6a164c) * $signed(16'hffff);
  assign T3565 = $signed(T3566) / $signed(22'h100000);
  assign T3566 = $signed(31'h2f05f637) * $signed(16'h0);
  assign T3567 = T2943[1'h0:1'h0];
  assign T3568 = T3577 ? twiddle4_3_83_imag : twiddle4_3_82_imag;
  assign twiddle4_3_82_imag = T3571 + T3569;
  assign T3569 = $signed(T3570) / $signed(22'h100000);
  assign T3570 = $signed(31'h2bd8692b) * $signed(16'hffff);
  assign T3571 = $signed(T3572) / $signed(22'h100000);
  assign T3572 = $signed(31'h2e9f291b) * $signed(16'h0);
  assign twiddle4_3_83_imag = T3575 + T3573;
  assign T3573 = $signed(T3574) / $signed(22'h100000);
  assign T3574 = $signed(31'h2c45c89f) * $signed(16'hffff);
  assign T3575 = $signed(T3576) / $signed(22'h100000);
  assign T3576 = $signed(31'h2e37592c) * $signed(16'h0);
  assign T3577 = T2943[1'h0:1'h0];
  assign T3578 = T2943[1'h1:1'h1];
  assign T3579 = T3600 ? T3590 : T3580;
  assign T3580 = T3589 ? twiddle4_3_85_imag : twiddle4_3_84_imag;
  assign twiddle4_3_84_imag = T3583 + T3581;
  assign T3581 = $signed(T3582) / $signed(22'h100000);
  assign T3582 = $signed(31'h2cb2324b) * $signed(16'hffff);
  assign T3583 = $signed(T3584) / $signed(22'h100000);
  assign T3584 = $signed(31'h2dce88a9) * $signed(16'h0);
  assign twiddle4_3_85_imag = T3587 + T3585;
  assign T3585 = $signed(T3586) / $signed(22'h100000);
  assign T3586 = $signed(31'h2d1da3d5) * $signed(16'hffff);
  assign T3587 = $signed(T3588) / $signed(22'h100000);
  assign T3588 = $signed(31'h2d64b9da) * $signed(16'h0);
  assign T3589 = T2943[1'h0:1'h0];
  assign T3590 = T3599 ? twiddle4_3_87_imag : twiddle4_3_86_imag;
  assign twiddle4_3_86_imag = T3593 + T3591;
  assign T3591 = $signed(T3592) / $signed(22'h100000);
  assign T3592 = $signed(31'h2d881ae7) * $signed(16'hffff);
  assign T3593 = $signed(T3594) / $signed(22'h100000);
  assign T3594 = $signed(31'h2cf9ef09) * $signed(16'h0);
  assign twiddle4_3_87_imag = T3597 + T3595;
  assign T3595 = $signed(T3596) / $signed(22'h100000);
  assign T3596 = $signed(31'h2df19533) * $signed(16'hffff);
  assign T3597 = $signed(T3598) / $signed(22'h100000);
  assign T3598 = $signed(31'h2c8e2a86) * $signed(16'h0);
  assign T3599 = T2943[1'h0:1'h0];
  assign T3600 = T2943[1'h1:1'h1];
  assign T3601 = T2943[2'h2:2'h2];
  assign T3602 = T3647 ? T3625 : T3603;
  assign T3603 = T3624 ? T3614 : T3604;
  assign T3604 = T3613 ? twiddle4_3_89_imag : twiddle4_3_88_imag;
  assign twiddle4_3_88_imag = T3607 + T3605;
  assign T3605 = $signed(T3606) / $signed(22'h100000);
  assign T3606 = $signed(31'h2e5a106f) * $signed(16'hffff);
  assign T3607 = $signed(T3608) / $signed(22'h100000);
  assign T3608 = $signed(31'h2c216eaa) * $signed(16'h0);
  assign twiddle4_3_89_imag = T3611 + T3609;
  assign T3609 = $signed(T3610) / $signed(22'h100000);
  assign T3610 = $signed(31'h2ec18a58) * $signed(16'hffff);
  assign T3611 = $signed(T3612) / $signed(22'h100000);
  assign T3612 = $signed(31'h2bb3bdce) * $signed(16'h0);
  assign T3613 = T2943[1'h0:1'h0];
  assign T3614 = T3623 ? twiddle4_3_91_imag : twiddle4_3_90_imag;
  assign twiddle4_3_90_imag = T3617 + T3615;
  assign T3615 = $signed(T3616) / $signed(22'h100000);
  assign T3616 = $signed(31'h2f2800ae) * $signed(16'hffff);
  assign T3617 = $signed(T3618) / $signed(22'h100000);
  assign T3618 = $signed(31'h2b451a54) * $signed(16'h0);
  assign twiddle4_3_91_imag = T3621 + T3619;
  assign T3619 = $signed(T3620) / $signed(22'h100000);
  assign T3620 = $signed(31'h2f8d7139) * $signed(16'hffff);
  assign T3621 = $signed(T3622) / $signed(22'h100000);
  assign T3622 = $signed(31'h2ad586a3) * $signed(16'h0);
  assign T3623 = T2943[1'h0:1'h0];
  assign T3624 = T2943[1'h1:1'h1];
  assign T3625 = T3646 ? T3636 : T3626;
  assign T3626 = T3635 ? twiddle4_3_93_imag : twiddle4_3_92_imag;
  assign twiddle4_3_92_imag = T3629 + T3627;
  assign T3627 = $signed(T3628) / $signed(22'h100000);
  assign T3628 = $signed(31'h2ff1d9c6) * $signed(16'hffff);
  assign T3629 = $signed(T3630) / $signed(22'h100000);
  assign T3630 = $signed(31'h2a650525) * $signed(16'h0);
  assign twiddle4_3_93_imag = T3633 + T3631;
  assign T3631 = $signed(T3632) / $signed(22'h100000);
  assign T3632 = $signed(31'h30553827) * $signed(16'hffff);
  assign T3633 = $signed(T3634) / $signed(22'h100000);
  assign T3634 = $signed(31'h29f3984b) * $signed(16'h0);
  assign T3635 = T2943[1'h0:1'h0];
  assign T3636 = T3645 ? twiddle4_3_95_imag : twiddle4_3_94_imag;
  assign twiddle4_3_94_imag = T3639 + T3637;
  assign T3637 = $signed(T3638) / $signed(22'h100000);
  assign T3638 = $signed(31'h30b78a35) * $signed(16'hffff);
  assign T3639 = $signed(T3640) / $signed(22'h100000);
  assign T3640 = $signed(31'h2981428b) * $signed(16'h0);
  assign twiddle4_3_95_imag = T3643 + T3641;
  assign T3641 = $signed(T3642) / $signed(22'h100000);
  assign T3642 = $signed(31'h3118cdce) * $signed(16'hffff);
  assign T3643 = $signed(T3644) / $signed(22'h100000);
  assign T3644 = $signed(31'h290e0660) * $signed(16'h0);
  assign T3645 = T2943[1'h0:1'h0];
  assign T3646 = T2943[1'h1:1'h1];
  assign T3647 = T2943[2'h2:2'h2];
  assign T3648 = T2943[2'h3:2'h3];
  assign T3649 = T2943[3'h4:3'h4];
  assign T3650 = T3867 ? T3745 : T3651;
  assign T3651 = T3744 ? T3698 : T3652;
  assign T3652 = T3697 ? T3675 : T3653;
  assign T3653 = T3674 ? T3664 : T3654;
  assign T3654 = T3663 ? twiddle4_3_97_imag : twiddle4_3_96_imag;
  assign twiddle4_3_96_imag = T3657 + T3655;
  assign T3655 = $signed(T3656) / $signed(22'h100000);
  assign T3656 = $signed(31'h317900d6) * $signed(16'hffff);
  assign T3657 = $signed(T3658) / $signed(22'h100000);
  assign T3658 = $signed(31'h2899e64a) * $signed(16'h0);
  assign twiddle4_3_97_imag = T3661 + T3659;
  assign T3659 = $signed(T3660) / $signed(22'h100000);
  assign T3660 = $signed(31'h31d82136) * $signed(16'hffff);
  assign T3661 = $signed(T3662) / $signed(22'h100000);
  assign T3662 = $signed(31'h2824e4cc) * $signed(16'h0);
  assign T3663 = T2943[1'h0:1'h0];
  assign T3664 = T3673 ? twiddle4_3_99_imag : twiddle4_3_98_imag;
  assign twiddle4_3_98_imag = T3667 + T3665;
  assign T3665 = $signed(T3666) / $signed(22'h100000);
  assign T3666 = $signed(31'h32362cdf) * $signed(16'hffff);
  assign T3667 = $signed(T3668) / $signed(22'h100000);
  assign T3668 = $signed(31'h27af0471) * $signed(16'h0);
  assign twiddle4_3_99_imag = T3671 + T3669;
  assign T3669 = $signed(T3670) / $signed(22'h100000);
  assign T3670 = $signed(31'h329321c7) * $signed(16'hffff);
  assign T3671 = $signed(T3672) / $signed(22'h100000);
  assign T3672 = $signed(31'h273847c7) * $signed(16'h0);
  assign T3673 = T2943[1'h0:1'h0];
  assign T3674 = T2943[1'h1:1'h1];
  assign T3675 = T3696 ? T3686 : T3676;
  assign T3676 = T3685 ? twiddle4_3_101_imag : twiddle4_3_100_imag;
  assign twiddle4_3_100_imag = T3679 + T3677;
  assign T3677 = $signed(T3678) / $signed(22'h100000);
  assign T3678 = $signed(31'h32eefde9) * $signed(16'hffff);
  assign T3679 = $signed(T3680) / $signed(22'h100000);
  assign T3680 = $signed(31'h26c0b162) * $signed(16'h0);
  assign twiddle4_3_101_imag = T3683 + T3681;
  assign T3681 = $signed(T3682) / $signed(22'h100000);
  assign T3682 = $signed(31'h3349bf48) * $signed(16'hffff);
  assign T3683 = $signed(T3684) / $signed(22'h100000);
  assign T3684 = $signed(31'h264843d8) * $signed(16'h0);
  assign T3685 = T2943[1'h0:1'h0];
  assign T3686 = T3695 ? twiddle4_3_103_imag : twiddle4_3_102_imag;
  assign twiddle4_3_102_imag = T3689 + T3687;
  assign T3687 = $signed(T3688) / $signed(22'h100000);
  assign T3688 = $signed(31'h33a363eb) * $signed(16'hffff);
  assign T3689 = $signed(T3690) / $signed(22'h100000);
  assign T3690 = $signed(31'h25cf01c7) * $signed(16'h0);
  assign twiddle4_3_103_imag = T3693 + T3691;
  assign T3691 = $signed(T3692) / $signed(22'h100000);
  assign T3692 = $signed(31'h33fbe9e2) * $signed(16'hffff);
  assign T3693 = $signed(T3694) / $signed(22'h100000);
  assign T3694 = $signed(31'h2554edd0) * $signed(16'h0);
  assign T3695 = T2943[1'h0:1'h0];
  assign T3696 = T2943[1'h1:1'h1];
  assign T3697 = T2943[2'h2:2'h2];
  assign T3698 = T3743 ? T3721 : T3699;
  assign T3699 = T3720 ? T3710 : T3700;
  assign T3700 = T3709 ? twiddle4_3_105_imag : twiddle4_3_104_imag;
  assign twiddle4_3_104_imag = T3703 + T3701;
  assign T3701 = $signed(T3702) / $signed(22'h100000);
  assign T3702 = $signed(31'h34534f40) * $signed(16'hffff);
  assign T3703 = $signed(T3704) / $signed(22'h100000);
  assign T3704 = $signed(31'h24da0a99) * $signed(16'h0);
  assign twiddle4_3_105_imag = T3707 + T3705;
  assign T3705 = $signed(T3706) / $signed(22'h100000);
  assign T3706 = $signed(31'h34a99221) * $signed(16'hffff);
  assign T3707 = $signed(T3708) / $signed(22'h100000);
  assign T3708 = $signed(31'h245e5acc) * $signed(16'h0);
  assign T3709 = T2943[1'h0:1'h0];
  assign T3710 = T3719 ? twiddle4_3_107_imag : twiddle4_3_106_imag;
  assign twiddle4_3_106_imag = T3713 + T3711;
  assign T3711 = $signed(T3712) / $signed(22'h100000);
  assign T3712 = $signed(31'h34feb0a5) * $signed(16'hffff);
  assign T3713 = $signed(T3714) / $signed(22'h100000);
  assign T3714 = $signed(31'h23e1e117) * $signed(16'h0);
  assign twiddle4_3_107_imag = T3717 + T3715;
  assign T3715 = $signed(T3716) / $signed(22'h100000);
  assign T3716 = $signed(31'h3552a8f4) * $signed(16'hffff);
  assign T3717 = $signed(T3718) / $signed(22'h100000);
  assign T3718 = $signed(31'h2364a02e) * $signed(16'h0);
  assign T3719 = T2943[1'h0:1'h0];
  assign T3720 = T2943[1'h1:1'h1];
  assign T3721 = T3742 ? T3732 : T3722;
  assign T3722 = T3731 ? twiddle4_3_109_imag : twiddle4_3_108_imag;
  assign twiddle4_3_108_imag = T3725 + T3723;
  assign T3723 = $signed(T3724) / $signed(22'h100000);
  assign T3724 = $signed(31'h35a5793c) * $signed(16'hffff);
  assign T3725 = $signed(T3726) / $signed(22'h100000);
  assign T3726 = $signed(31'h22e69ac7) * $signed(16'h0);
  assign twiddle4_3_109_imag = T3729 + T3727;
  assign T3727 = $signed(T3728) / $signed(22'h100000);
  assign T3728 = $signed(31'h35f71fb1) * $signed(16'hffff);
  assign T3729 = $signed(T3730) / $signed(22'h100000);
  assign T3730 = $signed(31'h2267d39f) * $signed(16'h0);
  assign T3731 = T2943[1'h0:1'h0];
  assign T3732 = T3741 ? twiddle4_3_111_imag : twiddle4_3_110_imag;
  assign twiddle4_3_110_imag = T3735 + T3733;
  assign T3733 = $signed(T3734) / $signed(22'h100000);
  assign T3734 = $signed(31'h36479a8e) * $signed(16'hffff);
  assign T3735 = $signed(T3736) / $signed(22'h100000);
  assign T3736 = $signed(31'h21e84d76) * $signed(16'h0);
  assign twiddle4_3_111_imag = T3739 + T3737;
  assign T3737 = $signed(T3738) / $signed(22'h100000);
  assign T3738 = $signed(31'h3696e813) * $signed(16'hffff);
  assign T3739 = $signed(T3740) / $signed(22'h100000);
  assign T3740 = $signed(31'h21680b0f) * $signed(16'h0);
  assign T3741 = T2943[1'h0:1'h0];
  assign T3742 = T2943[1'h1:1'h1];
  assign T3743 = T2943[2'h2:2'h2];
  assign T3744 = T2943[2'h3:2'h3];
  assign T3745 = T3866 ? T3804 : T3746;
  assign T3746 = T3803 ? T3773 : T3747;
  assign T3747 = T3772 ? T3758 : T3748;
  assign T3748 = T3757 ? twiddle4_3_113_imag : twiddle4_3_112_imag;
  assign twiddle4_3_112_imag = T3751 + T3749;
  assign T3749 = $signed(T3750) / $signed(22'h100000);
  assign T3750 = $signed(31'h36e5068a) * $signed(16'hffff);
  assign T3751 = $signed(T3752) / $signed(22'h100000);
  assign T3752 = $signed(31'h20e70f32) * $signed(16'h0);
  assign twiddle4_3_113_imag = T3755 + T3753;
  assign T3753 = $signed(T3754) / $signed(22'h100000);
  assign T3754 = $signed(31'h3731f43f) * $signed(16'hffff);
  assign T3755 = $signed(T3756) / $signed(22'h100000);
  assign T3756 = $signed(31'h20655cab) * $signed(16'h0);
  assign T3757 = T2943[1'h0:1'h0];
  assign T3758 = T3771 ? twiddle4_3_115_imag : twiddle4_3_114_imag;
  assign twiddle4_3_114_imag = T3761 + T3759;
  assign T3759 = $signed(T3760) / $signed(22'h100000);
  assign T3760 = $signed(31'h377daf89) * $signed(16'hffff);
  assign T3761 = {T3764, T3762};
  assign T3762 = $signed(T3763) / $signed(22'h100000);
  assign T3763 = $signed(30'h1fe2f64b) * $signed(16'h0);
  assign T3764 = T3762[6'h2d:6'h2d];
  assign twiddle4_3_115_imag = T3767 + T3765;
  assign T3765 = $signed(T3766) / $signed(22'h100000);
  assign T3766 = $signed(31'h37c836c2) * $signed(16'hffff);
  assign T3767 = {T3770, T3768};
  assign T3768 = $signed(T3769) / $signed(22'h100000);
  assign T3769 = $signed(30'h1f5fdee6) * $signed(16'h0);
  assign T3770 = T3768[6'h2d:6'h2d];
  assign T3771 = T2943[1'h0:1'h0];
  assign T3772 = T2943[1'h1:1'h1];
  assign T3773 = T3802 ? T3788 : T3774;
  assign T3774 = T3787 ? twiddle4_3_117_imag : twiddle4_3_116_imag;
  assign twiddle4_3_116_imag = T3777 + T3775;
  assign T3775 = $signed(T3776) / $signed(22'h100000);
  assign T3776 = $signed(31'h3811884c) * $signed(16'hffff);
  assign T3777 = {T3780, T3778};
  assign T3778 = $signed(T3779) / $signed(22'h100000);
  assign T3779 = $signed(30'h1edc1952) * $signed(16'h0);
  assign T3780 = T3778[6'h2d:6'h2d];
  assign twiddle4_3_117_imag = T3783 + T3781;
  assign T3781 = $signed(T3782) / $signed(22'h100000);
  assign T3782 = $signed(31'h3859a292) * $signed(16'hffff);
  assign T3783 = {T3786, T3784};
  assign T3784 = $signed(T3785) / $signed(22'h100000);
  assign T3785 = $signed(30'h1e57a86d) * $signed(16'h0);
  assign T3786 = T3784[6'h2d:6'h2d];
  assign T3787 = T2943[1'h0:1'h0];
  assign T3788 = T3801 ? twiddle4_3_119_imag : twiddle4_3_118_imag;
  assign twiddle4_3_118_imag = T3791 + T3789;
  assign T3789 = $signed(T3790) / $signed(22'h100000);
  assign T3790 = $signed(31'h38a08402) * $signed(16'hffff);
  assign T3791 = {T3794, T3792};
  assign T3792 = $signed(T3793) / $signed(22'h100000);
  assign T3793 = $signed(30'h1dd28f14) * $signed(16'h0);
  assign T3794 = T3792[6'h2d:6'h2d];
  assign twiddle4_3_119_imag = T3797 + T3795;
  assign T3795 = $signed(T3796) / $signed(22'h100000);
  assign T3796 = $signed(31'h38e62b13) * $signed(16'hffff);
  assign T3797 = {T3800, T3798};
  assign T3798 = $signed(T3799) / $signed(22'h100000);
  assign T3799 = $signed(30'h1d4cd02b) * $signed(16'h0);
  assign T3800 = T3798[6'h2d:6'h2d];
  assign T3801 = T2943[1'h0:1'h0];
  assign T3802 = T2943[1'h1:1'h1];
  assign T3803 = T2943[2'h2:2'h2];
  assign T3804 = T3865 ? T3835 : T3805;
  assign T3805 = T3834 ? T3820 : T3806;
  assign T3806 = T3819 ? twiddle4_3_121_imag : twiddle4_3_120_imag;
  assign twiddle4_3_120_imag = T3809 + T3807;
  assign T3807 = $signed(T3808) / $signed(22'h100000);
  assign T3808 = $signed(31'h392a9642) * $signed(16'hffff);
  assign T3809 = {T3812, T3810};
  assign T3810 = $signed(T3811) / $signed(22'h100000);
  assign T3811 = $signed(30'h1cc66e99) * $signed(16'h0);
  assign T3812 = T3810[6'h2d:6'h2d];
  assign twiddle4_3_121_imag = T3815 + T3813;
  assign T3813 = $signed(T3814) / $signed(22'h100000);
  assign T3814 = $signed(31'h396dc414) * $signed(16'hffff);
  assign T3815 = {T3818, T3816};
  assign T3816 = $signed(T3817) / $signed(22'h100000);
  assign T3817 = $signed(30'h1c3f6d47) * $signed(16'h0);
  assign T3818 = T3816[6'h2d:6'h2d];
  assign T3819 = T2943[1'h0:1'h0];
  assign T3820 = T3833 ? twiddle4_3_123_imag : twiddle4_3_122_imag;
  assign twiddle4_3_122_imag = T3823 + T3821;
  assign T3821 = $signed(T3822) / $signed(22'h100000);
  assign T3822 = $signed(31'h39afb313) * $signed(16'hffff);
  assign T3823 = {T3826, T3824};
  assign T3824 = $signed(T3825) / $signed(22'h100000);
  assign T3825 = $signed(30'h1bb7cf23) * $signed(16'h0);
  assign T3826 = T3824[6'h2d:6'h2d];
  assign twiddle4_3_123_imag = T3829 + T3827;
  assign T3827 = $signed(T3828) / $signed(22'h100000);
  assign T3828 = $signed(31'h39f061d1) * $signed(16'hffff);
  assign T3829 = {T3832, T3830};
  assign T3830 = $signed(T3831) / $signed(22'h100000);
  assign T3831 = $signed(30'h1b2f971d) * $signed(16'h0);
  assign T3832 = T3830[6'h2d:6'h2d];
  assign T3833 = T2943[1'h0:1'h0];
  assign T3834 = T2943[1'h1:1'h1];
  assign T3835 = T3864 ? T3850 : T3836;
  assign T3836 = T3849 ? twiddle4_3_125_imag : twiddle4_3_124_imag;
  assign twiddle4_3_124_imag = T3839 + T3837;
  assign T3837 = $signed(T3838) / $signed(22'h100000);
  assign T3838 = $signed(31'h3a2fcee8) * $signed(16'hffff);
  assign T3839 = {T3842, T3840};
  assign T3840 = $signed(T3841) / $signed(22'h100000);
  assign T3841 = $signed(30'h1aa6c82b) * $signed(16'h0);
  assign T3842 = T3840[6'h2d:6'h2d];
  assign twiddle4_3_125_imag = T3845 + T3843;
  assign T3843 = $signed(T3844) / $signed(22'h100000);
  assign T3844 = $signed(31'h3a6df8f7) * $signed(16'hffff);
  assign T3845 = {T3848, T3846};
  assign T3846 = $signed(T3847) / $signed(22'h100000);
  assign T3847 = $signed(30'h1a1d6543) * $signed(16'h0);
  assign T3848 = T3846[6'h2d:6'h2d];
  assign T3849 = T2943[1'h0:1'h0];
  assign T3850 = T3863 ? twiddle4_3_127_imag : twiddle4_3_126_imag;
  assign twiddle4_3_126_imag = T3853 + T3851;
  assign T3851 = $signed(T3852) / $signed(22'h100000);
  assign T3852 = $signed(31'h3aaadea5) * $signed(16'hffff);
  assign T3853 = {T3856, T3854};
  assign T3854 = $signed(T3855) / $signed(22'h100000);
  assign T3855 = $signed(30'h19937161) * $signed(16'h0);
  assign T3856 = T3854[6'h2d:6'h2d];
  assign twiddle4_3_127_imag = T3859 + T3857;
  assign T3857 = $signed(T3858) / $signed(22'h100000);
  assign T3858 = $signed(31'h3ae67ea1) * $signed(16'hffff);
  assign T3859 = {T3862, T3860};
  assign T3860 = $signed(T3861) / $signed(22'h100000);
  assign T3861 = $signed(30'h1908ef81) * $signed(16'h0);
  assign T3862 = T3860[6'h2d:6'h2d];
  assign T3863 = T2943[1'h0:1'h0];
  assign T3864 = T2943[1'h1:1'h1];
  assign T3865 = T2943[2'h2:2'h2];
  assign T3866 = T2943[2'h3:2'h3];
  assign T3867 = T2943[3'h4:3'h4];
  assign T3868 = T2943[3'h5:3'h5];
  assign T3869 = T3459[6'h2e:6'h2e];
  assign T3870 = T2943[3'h6:3'h6];
  assign T3871 = {T4893, T3872};
  assign T3872 = T4892 ? T4431 : T3873;
  assign T3873 = T4430 ? T4144 : T3874;
  assign T3874 = T4143 ? T4001 : T3875;
  assign T3875 = T4000 ? T3938 : T3876;
  assign T3876 = T3937 ? T3907 : T3877;
  assign T3877 = T3906 ? T3892 : T3878;
  assign T3878 = T3891 ? twiddle4_3_129_imag : twiddle4_3_128_imag;
  assign twiddle4_3_128_imag = T3881 + T3879;
  assign T3879 = $signed(T3880) / $signed(22'h100000);
  assign T3880 = $signed(31'h3b20d79e) * $signed(16'hffff);
  assign T3881 = {T3884, T3882};
  assign T3882 = $signed(T3883) / $signed(22'h100000);
  assign T3883 = $signed(30'h187de2a6) * $signed(16'h0);
  assign T3884 = T3882[6'h2d:6'h2d];
  assign twiddle4_3_129_imag = T3887 + T3885;
  assign T3885 = $signed(T3886) / $signed(22'h100000);
  assign T3886 = $signed(31'h3b59e859) * $signed(16'hffff);
  assign T3887 = {T3890, T3888};
  assign T3888 = $signed(T3889) / $signed(22'h100000);
  assign T3889 = $signed(30'h17f24dd3) * $signed(16'h0);
  assign T3890 = T3888[6'h2d:6'h2d];
  assign T3891 = T2943[1'h0:1'h0];
  assign T3892 = T3905 ? twiddle4_3_131_imag : twiddle4_3_130_imag;
  assign twiddle4_3_130_imag = T3895 + T3893;
  assign T3893 = $signed(T3894) / $signed(22'h100000);
  assign T3894 = $signed(31'h3b91af96) * $signed(16'hffff);
  assign T3895 = {T3898, T3896};
  assign T3896 = $signed(T3897) / $signed(22'h100000);
  assign T3897 = $signed(30'h1766340f) * $signed(16'h0);
  assign T3898 = T3896[6'h2d:6'h2d];
  assign twiddle4_3_131_imag = T3901 + T3899;
  assign T3899 = $signed(T3900) / $signed(22'h100000);
  assign T3900 = $signed(31'h3bc82c1e) * $signed(16'hffff);
  assign T3901 = {T3904, T3902};
  assign T3902 = $signed(T3903) / $signed(22'h100000);
  assign T3903 = $signed(30'h16d99863) * $signed(16'h0);
  assign T3904 = T3902[6'h2d:6'h2d];
  assign T3905 = T2943[1'h0:1'h0];
  assign T3906 = T2943[1'h1:1'h1];
  assign T3907 = T3936 ? T3922 : T3908;
  assign T3908 = T3921 ? twiddle4_3_133_imag : twiddle4_3_132_imag;
  assign twiddle4_3_132_imag = T3911 + T3909;
  assign T3909 = $signed(T3910) / $signed(22'h100000);
  assign T3910 = $signed(31'h3bfd5cc4) * $signed(16'hffff);
  assign T3911 = {T3914, T3912};
  assign T3912 = $signed(T3913) / $signed(22'h100000);
  assign T3913 = $signed(30'h164c7ddd) * $signed(16'h0);
  assign T3914 = T3912[6'h2d:6'h2d];
  assign twiddle4_3_133_imag = T3917 + T3915;
  assign T3915 = $signed(T3916) / $signed(22'h100000);
  assign T3916 = $signed(31'h3c31405f) * $signed(16'hffff);
  assign T3917 = {T3920, T3918};
  assign T3918 = $signed(T3919) / $signed(22'h100000);
  assign T3919 = $signed(30'h15bee78b) * $signed(16'h0);
  assign T3920 = T3918[6'h2d:6'h2d];
  assign T3921 = T2943[1'h0:1'h0];
  assign T3922 = T3935 ? twiddle4_3_135_imag : twiddle4_3_134_imag;
  assign twiddle4_3_134_imag = T3925 + T3923;
  assign T3923 = $signed(T3924) / $signed(22'h100000);
  assign T3924 = $signed(31'h3c63d5d0) * $signed(16'hffff);
  assign T3925 = {T3928, T3926};
  assign T3926 = $signed(T3927) / $signed(22'h100000);
  assign T3927 = $signed(30'h1530d880) * $signed(16'h0);
  assign T3928 = T3926[6'h2d:6'h2d];
  assign twiddle4_3_135_imag = T3931 + T3929;
  assign T3929 = $signed(T3930) / $signed(22'h100000);
  assign T3930 = $signed(31'h3c951bff) * $signed(16'hffff);
  assign T3931 = {T3934, T3932};
  assign T3932 = $signed(T3933) / $signed(22'h100000);
  assign T3933 = $signed(30'h14a253d1) * $signed(16'h0);
  assign T3934 = T3932[6'h2d:6'h2d];
  assign T3935 = T2943[1'h0:1'h0];
  assign T3936 = T2943[1'h1:1'h1];
  assign T3937 = T2943[2'h2:2'h2];
  assign T3938 = T3999 ? T3969 : T3939;
  assign T3939 = T3968 ? T3954 : T3940;
  assign T3940 = T3953 ? twiddle4_3_137_imag : twiddle4_3_136_imag;
  assign twiddle4_3_136_imag = T3943 + T3941;
  assign T3941 = $signed(T3942) / $signed(22'h100000);
  assign T3942 = $signed(31'h3cc511d8) * $signed(16'hffff);
  assign T3943 = {T3946, T3944};
  assign T3944 = $signed(T3945) / $signed(22'h100000);
  assign T3945 = $signed(30'h14135c94) * $signed(16'h0);
  assign T3946 = T3944[6'h2d:6'h2d];
  assign twiddle4_3_137_imag = T3949 + T3947;
  assign T3947 = $signed(T3948) / $signed(22'h100000);
  assign T3948 = $signed(31'h3cf3b653) * $signed(16'hffff);
  assign T3949 = {T3952, T3950};
  assign T3950 = $signed(T3951) / $signed(22'h100000);
  assign T3951 = $signed(30'h1383f5e3) * $signed(16'h0);
  assign T3952 = T3950[6'h2d:6'h2d];
  assign T3953 = T2943[1'h0:1'h0];
  assign T3954 = T3967 ? twiddle4_3_139_imag : twiddle4_3_138_imag;
  assign twiddle4_3_138_imag = T3957 + T3955;
  assign T3955 = $signed(T3956) / $signed(22'h100000);
  assign T3956 = $signed(31'h3d21086c) * $signed(16'hffff);
  assign T3957 = {T3960, T3958};
  assign T3958 = $signed(T3959) / $signed(22'h100000);
  assign T3959 = $signed(30'h12f422da) * $signed(16'h0);
  assign T3960 = T3958[6'h2d:6'h2d];
  assign twiddle4_3_139_imag = T3963 + T3961;
  assign T3961 = $signed(T3962) / $signed(22'h100000);
  assign T3962 = $signed(31'h3d4d0727) * $signed(16'hffff);
  assign T3963 = {T3966, T3964};
  assign T3964 = $signed(T3965) / $signed(22'h100000);
  assign T3965 = $signed(30'h1263e699) * $signed(16'h0);
  assign T3966 = T3964[6'h2d:6'h2d];
  assign T3967 = T2943[1'h0:1'h0];
  assign T3968 = T2943[1'h1:1'h1];
  assign T3969 = T3998 ? T3984 : T3970;
  assign T3970 = T3983 ? twiddle4_3_141_imag : twiddle4_3_140_imag;
  assign twiddle4_3_140_imag = T3973 + T3971;
  assign T3971 = $signed(T3972) / $signed(22'h100000);
  assign T3972 = $signed(31'h3d77b191) * $signed(16'hffff);
  assign T3973 = {T3976, T3974};
  assign T3974 = $signed(T3975) / $signed(22'h100000);
  assign T3975 = $signed(30'h11d3443f) * $signed(16'h0);
  assign T3976 = T3974[6'h2d:6'h2d];
  assign twiddle4_3_141_imag = T3979 + T3977;
  assign T3977 = $signed(T3978) / $signed(22'h100000);
  assign T3978 = $signed(31'h3da106bd) * $signed(16'hffff);
  assign T3979 = {T3982, T3980};
  assign T3980 = $signed(T3981) / $signed(22'h100000);
  assign T3981 = $signed(30'h11423eef) * $signed(16'h0);
  assign T3982 = T3980[6'h2d:6'h2d];
  assign T3983 = T2943[1'h0:1'h0];
  assign T3984 = T3997 ? twiddle4_3_143_imag : twiddle4_3_142_imag;
  assign twiddle4_3_142_imag = T3987 + T3985;
  assign T3985 = $signed(T3986) / $signed(22'h100000);
  assign T3986 = $signed(31'h3dc905c4) * $signed(16'hffff);
  assign T3987 = {T3990, T3988};
  assign T3988 = $signed(T3989) / $signed(22'h100000);
  assign T3989 = $signed(30'h10b0d9cf) * $signed(16'h0);
  assign T3990 = T3988[6'h2d:6'h2d];
  assign twiddle4_3_143_imag = T3993 + T3991;
  assign T3991 = $signed(T3992) / $signed(22'h100000);
  assign T3992 = $signed(31'h3defadca) * $signed(16'hffff);
  assign T3993 = {T3996, T3994};
  assign T3994 = $signed(T3995) / $signed(22'h100000);
  assign T3995 = $signed(30'h101f1806) * $signed(16'h0);
  assign T3996 = T3994[6'h2d:6'h2d];
  assign T3997 = T2943[1'h0:1'h0];
  assign T3998 = T2943[1'h1:1'h1];
  assign T3999 = T2943[2'h2:2'h2];
  assign T4000 = T2943[2'h3:2'h3];
  assign T4001 = T4142 ? T4072 : T4002;
  assign T4002 = T4071 ? T4037 : T4003;
  assign T4003 = T4036 ? T4020 : T4004;
  assign T4004 = T4019 ? twiddle4_3_145_imag : twiddle4_3_144_imag;
  assign twiddle4_3_144_imag = T4007 + T4005;
  assign T4005 = $signed(T4006) / $signed(22'h100000);
  assign T4006 = $signed(31'h3e14fdf7) * $signed(16'hffff);
  assign T4007 = {T4010, T4008};
  assign T4008 = $signed(T4009) / $signed(22'h100000);
  assign T4009 = $signed(29'hf8cfcbd) * $signed(16'h0);
  assign T4010 = T4011 ? 2'h3 : 2'h0;
  assign T4011 = T4008[6'h2c:6'h2c];
  assign twiddle4_3_145_imag = T4014 + T4012;
  assign T4012 = $signed(T4013) / $signed(22'h100000);
  assign T4013 = $signed(31'h3e38f57c) * $signed(16'hffff);
  assign T4014 = {T4017, T4015};
  assign T4015 = $signed(T4016) / $signed(22'h100000);
  assign T4016 = $signed(29'hefa8b1f) * $signed(16'h0);
  assign T4017 = T4018 ? 2'h3 : 2'h0;
  assign T4018 = T4015[6'h2c:6'h2c];
  assign T4019 = T2943[1'h0:1'h0];
  assign T4020 = T4035 ? twiddle4_3_147_imag : twiddle4_3_146_imag;
  assign twiddle4_3_146_imag = T4023 + T4021;
  assign T4021 = $signed(T4022) / $signed(22'h100000);
  assign T4022 = $signed(31'h3e5b9392) * $signed(16'hffff);
  assign T4023 = {T4026, T4024};
  assign T4024 = $signed(T4025) / $signed(22'h100000);
  assign T4025 = $signed(29'he67c659) * $signed(16'h0);
  assign T4026 = T4027 ? 2'h3 : 2'h0;
  assign T4027 = T4024[6'h2c:6'h2c];
  assign twiddle4_3_147_imag = T4030 + T4028;
  assign T4028 = $signed(T4029) / $signed(22'h100000);
  assign T4029 = $signed(31'h3e7cd778) * $signed(16'hffff);
  assign T4030 = {T4033, T4031};
  assign T4031 = $signed(T4032) / $signed(22'h100000);
  assign T4032 = $signed(29'hdd4b19a) * $signed(16'h0);
  assign T4033 = T4034 ? 2'h3 : 2'h0;
  assign T4034 = T4031[6'h2c:6'h2c];
  assign T4035 = T2943[1'h0:1'h0];
  assign T4036 = T2943[1'h1:1'h1];
  assign T4037 = T4070 ? T4054 : T4038;
  assign T4038 = T4053 ? twiddle4_3_149_imag : twiddle4_3_148_imag;
  assign twiddle4_3_148_imag = T4041 + T4039;
  assign T4039 = $signed(T4040) / $signed(22'h100000);
  assign T4040 = $signed(31'h3e9cc076) * $signed(16'hffff);
  assign T4041 = {T4044, T4042};
  assign T4042 = $signed(T4043) / $signed(22'h100000);
  assign T4043 = $signed(29'hd415012) * $signed(16'h0);
  assign T4044 = T4045 ? 2'h3 : 2'h0;
  assign T4045 = T4042[6'h2c:6'h2c];
  assign twiddle4_3_149_imag = T4048 + T4046;
  assign T4046 = $signed(T4047) / $signed(22'h100000);
  assign T4047 = $signed(31'h3ebb4dda) * $signed(16'hffff);
  assign T4048 = {T4051, T4049};
  assign T4049 = $signed(T4050) / $signed(22'h100000);
  assign T4050 = $signed(29'hcada4f4) * $signed(16'h0);
  assign T4051 = T4052 ? 2'h3 : 2'h0;
  assign T4052 = T4049[6'h2c:6'h2c];
  assign T4053 = T2943[1'h0:1'h0];
  assign T4054 = T4069 ? twiddle4_3_151_imag : twiddle4_3_150_imag;
  assign twiddle4_3_150_imag = T4057 + T4055;
  assign T4055 = $signed(T4056) / $signed(22'h100000);
  assign T4056 = $signed(31'h3ed87efb) * $signed(16'hffff);
  assign T4057 = {T4060, T4058};
  assign T4058 = $signed(T4059) / $signed(22'h100000);
  assign T4059 = $signed(29'hc19b374) * $signed(16'h0);
  assign T4060 = T4061 ? 2'h3 : 2'h0;
  assign T4061 = T4058[6'h2c:6'h2c];
  assign twiddle4_3_151_imag = T4064 + T4062;
  assign T4062 = $signed(T4063) / $signed(22'h100000);
  assign T4063 = $signed(31'h3ef45338) * $signed(16'hffff);
  assign T4064 = {T4067, T4065};
  assign T4065 = $signed(T4066) / $signed(22'h100000);
  assign T4066 = $signed(29'hb857ec6) * $signed(16'h0);
  assign T4067 = T4068 ? 2'h3 : 2'h0;
  assign T4068 = T4065[6'h2c:6'h2c];
  assign T4069 = T2943[1'h0:1'h0];
  assign T4070 = T2943[1'h1:1'h1];
  assign T4071 = T2943[2'h2:2'h2];
  assign T4072 = T4141 ? T4107 : T4073;
  assign T4073 = T4106 ? T4090 : T4074;
  assign T4074 = T4089 ? twiddle4_3_153_imag : twiddle4_3_152_imag;
  assign twiddle4_3_152_imag = T4077 + T4075;
  assign T4075 = $signed(T4076) / $signed(22'h100000);
  assign T4076 = $signed(31'h3f0ec9f4) * $signed(16'hffff);
  assign T4077 = {T4080, T4078};
  assign T4078 = $signed(T4079) / $signed(22'h100000);
  assign T4079 = $signed(29'haf10a22) * $signed(16'h0);
  assign T4080 = T4081 ? 2'h3 : 2'h0;
  assign T4081 = T4078[6'h2c:6'h2c];
  assign twiddle4_3_153_imag = T4084 + T4082;
  assign T4082 = $signed(T4083) / $signed(22'h100000);
  assign T4083 = $signed(31'h3f27e29f) * $signed(16'hffff);
  assign T4084 = {T4087, T4085};
  assign T4085 = $signed(T4086) / $signed(22'h100000);
  assign T4086 = $signed(29'ha5c58bf) * $signed(16'h0);
  assign T4087 = T4088 ? 2'h3 : 2'h0;
  assign T4088 = T4085[6'h2c:6'h2c];
  assign T4089 = T2943[1'h0:1'h0];
  assign T4090 = T4105 ? twiddle4_3_155_imag : twiddle4_3_154_imag;
  assign twiddle4_3_154_imag = T4093 + T4091;
  assign T4091 = $signed(T4092) / $signed(22'h100000);
  assign T4092 = $signed(31'h3f3f9cab) * $signed(16'hffff);
  assign T4093 = {T4096, T4094};
  assign T4094 = $signed(T4095) / $signed(22'h100000);
  assign T4095 = $signed(29'h9c76dd8) * $signed(16'h0);
  assign T4096 = T4097 ? 2'h3 : 2'h0;
  assign T4097 = T4094[6'h2c:6'h2c];
  assign twiddle4_3_155_imag = T4100 + T4098;
  assign T4098 = $signed(T4099) / $signed(22'h100000);
  assign T4099 = $signed(31'h3f55f796) * $signed(16'hffff);
  assign T4100 = {T4103, T4101};
  assign T4101 = $signed(T4102) / $signed(22'h100000);
  assign T4102 = $signed(29'h9324ca6) * $signed(16'h0);
  assign T4103 = T4104 ? 2'h3 : 2'h0;
  assign T4104 = T4101[6'h2c:6'h2c];
  assign T4105 = T2943[1'h0:1'h0];
  assign T4106 = T2943[1'h1:1'h1];
  assign T4107 = T4140 ? T4124 : T4108;
  assign T4108 = T4123 ? twiddle4_3_157_imag : twiddle4_3_156_imag;
  assign twiddle4_3_156_imag = T4111 + T4109;
  assign T4109 = $signed(T4110) / $signed(22'h100000);
  assign T4110 = $signed(31'h3f6af2e3) * $signed(16'hffff);
  assign T4111 = {T4114, T4112};
  assign T4112 = $signed(T4113) / $signed(22'h100000);
  assign T4113 = $signed(29'h89cf867) * $signed(16'h0);
  assign T4114 = T4115 ? 2'h3 : 2'h0;
  assign T4115 = T4112[6'h2c:6'h2c];
  assign twiddle4_3_157_imag = T4118 + T4116;
  assign T4116 = $signed(T4117) / $signed(22'h100000);
  assign T4117 = $signed(31'h3f7e8e1e) * $signed(16'hffff);
  assign T4118 = {T4121, T4119};
  assign T4119 = $signed(T4120) / $signed(22'h100000);
  assign T4120 = $signed(29'h8077456) * $signed(16'h0);
  assign T4121 = T4122 ? 2'h3 : 2'h0;
  assign T4122 = T4119[6'h2c:6'h2c];
  assign T4123 = T2943[1'h0:1'h0];
  assign T4124 = T4139 ? twiddle4_3_159_imag : twiddle4_3_158_imag;
  assign twiddle4_3_158_imag = T4127 + T4125;
  assign T4125 = $signed(T4126) / $signed(22'h100000);
  assign T4126 = $signed(31'h3f90c8d9) * $signed(16'hffff);
  assign T4127 = {T4130, T4128};
  assign T4128 = $signed(T4129) / $signed(22'h100000);
  assign T4129 = $signed(28'h771c3b2) * $signed(16'h0);
  assign T4130 = T4131 ? 3'h7 : 3'h0;
  assign T4131 = T4128[6'h2b:6'h2b];
  assign twiddle4_3_159_imag = T4134 + T4132;
  assign T4132 = $signed(T4133) / $signed(22'h100000);
  assign T4133 = $signed(31'h3fa1a2b1) * $signed(16'hffff);
  assign T4134 = {T4137, T4135};
  assign T4135 = $signed(T4136) / $signed(22'h100000);
  assign T4136 = $signed(28'h6dbe9bb) * $signed(16'h0);
  assign T4137 = T4138 ? 3'h7 : 3'h0;
  assign T4138 = T4135[6'h2b:6'h2b];
  assign T4139 = T2943[1'h0:1'h0];
  assign T4140 = T2943[1'h1:1'h1];
  assign T4141 = T2943[2'h2:2'h2];
  assign T4142 = T2943[2'h3:2'h3];
  assign T4143 = T2943[3'h4:3'h4];
  assign T4144 = T4429 ? T4287 : T4145;
  assign T4145 = T4286 ? T4216 : T4146;
  assign T4146 = T4215 ? T4181 : T4147;
  assign T4147 = T4180 ? T4164 : T4148;
  assign T4148 = T4163 ? twiddle4_3_161_imag : twiddle4_3_160_imag;
  assign twiddle4_3_160_imag = T4151 + T4149;
  assign T4149 = $signed(T4150) / $signed(22'h100000);
  assign T4150 = $signed(31'h3fb11b47) * $signed(16'hffff);
  assign T4151 = {T4154, T4152};
  assign T4152 = $signed(T4153) / $signed(22'h100000);
  assign T4153 = $signed(28'h645e9af) * $signed(16'h0);
  assign T4154 = T4155 ? 3'h7 : 3'h0;
  assign T4155 = T4152[6'h2b:6'h2b];
  assign twiddle4_3_161_imag = T4158 + T4156;
  assign T4156 = $signed(T4157) / $signed(22'h100000);
  assign T4157 = $signed(31'h3fbf3245) * $signed(16'hffff);
  assign T4158 = {T4161, T4159};
  assign T4159 = $signed(T4160) / $signed(22'h100000);
  assign T4160 = $signed(28'h5afc6cf) * $signed(16'h0);
  assign T4161 = T4162 ? 3'h7 : 3'h0;
  assign T4162 = T4159[6'h2b:6'h2b];
  assign T4163 = T2943[1'h0:1'h0];
  assign T4164 = T4179 ? twiddle4_3_163_imag : twiddle4_3_162_imag;
  assign twiddle4_3_162_imag = T4167 + T4165;
  assign T4165 = $signed(T4166) / $signed(22'h100000);
  assign T4166 = $signed(31'h3fcbe75e) * $signed(16'hffff);
  assign T4167 = {T4170, T4168};
  assign T4168 = $signed(T4169) / $signed(22'h100000);
  assign T4169 = $signed(28'h519845e) * $signed(16'h0);
  assign T4170 = T4171 ? 3'h7 : 3'h0;
  assign T4171 = T4168[6'h2b:6'h2b];
  assign twiddle4_3_163_imag = T4174 + T4172;
  assign T4172 = $signed(T4173) / $signed(22'h100000);
  assign T4173 = $signed(31'h3fd73a4a) * $signed(16'hffff);
  assign T4174 = {T4177, T4175};
  assign T4175 = $signed(T4176) / $signed(22'h100000);
  assign T4176 = $signed(28'h483259d) * $signed(16'h0);
  assign T4177 = T4178 ? 3'h7 : 3'h0;
  assign T4178 = T4175[6'h2b:6'h2b];
  assign T4179 = T2943[1'h0:1'h0];
  assign T4180 = T2943[1'h1:1'h1];
  assign T4181 = T4214 ? T4198 : T4182;
  assign T4182 = T4197 ? twiddle4_3_165_imag : twiddle4_3_164_imag;
  assign twiddle4_3_164_imag = T4185 + T4183;
  assign T4183 = $signed(T4184) / $signed(22'h100000);
  assign T4184 = $signed(31'h3fe12acb) * $signed(16'hffff);
  assign T4185 = {T4188, T4186};
  assign T4186 = $signed(T4187) / $signed(22'h100000);
  assign T4187 = $signed(27'h3ecadcf) * $signed(16'h0);
  assign T4188 = T4189 ? 4'hf : 4'h0;
  assign T4189 = T4186[6'h2a:6'h2a];
  assign twiddle4_3_165_imag = T4192 + T4190;
  assign T4190 = $signed(T4191) / $signed(22'h100000);
  assign T4191 = $signed(31'h3fe9b8a9) * $signed(16'hffff);
  assign T4192 = {T4195, T4193};
  assign T4193 = $signed(T4194) / $signed(22'h100000);
  assign T4194 = $signed(27'h3562037) * $signed(16'h0);
  assign T4195 = T4196 ? 4'hf : 4'h0;
  assign T4196 = T4193[6'h2a:6'h2a];
  assign T4197 = T2943[1'h0:1'h0];
  assign T4198 = T4213 ? twiddle4_3_167_imag : twiddle4_3_166_imag;
  assign twiddle4_3_166_imag = T4201 + T4199;
  assign T4199 = $signed(T4200) / $signed(22'h100000);
  assign T4200 = $signed(31'h3ff0e3b5) * $signed(16'hffff);
  assign T4201 = {T4204, T4202};
  assign T4202 = $signed(T4203) / $signed(22'h100000);
  assign T4203 = $signed(27'h2bf801a) * $signed(16'h0);
  assign T4204 = T4205 ? 4'hf : 4'h0;
  assign T4205 = T4202[6'h2a:6'h2a];
  assign twiddle4_3_167_imag = T4208 + T4206;
  assign T4206 = $signed(T4207) / $signed(22'h100000);
  assign T4207 = $signed(31'h3ff6abc8) * $signed(16'hffff);
  assign T4208 = {T4211, T4209};
  assign T4209 = $signed(T4210) / $signed(22'h100000);
  assign T4210 = $signed(27'h228d0bb) * $signed(16'h0);
  assign T4211 = T4212 ? 4'hf : 4'h0;
  assign T4212 = T4209[6'h2a:6'h2a];
  assign T4213 = T2943[1'h0:1'h0];
  assign T4214 = T2943[1'h1:1'h1];
  assign T4215 = T2943[2'h2:2'h2];
  assign T4216 = T4285 ? T4251 : T4217;
  assign T4217 = T4250 ? T4234 : T4218;
  assign T4218 = T4233 ? twiddle4_3_169_imag : twiddle4_3_168_imag;
  assign twiddle4_3_168_imag = T4221 + T4219;
  assign T4219 = $signed(T4220) / $signed(22'h100000);
  assign T4220 = $signed(31'h3ffb10c1) * $signed(16'hffff);
  assign T4221 = {T4224, T4222};
  assign T4222 = $signed(T4223) / $signed(22'h100000);
  assign T4223 = $signed(26'h192155f) * $signed(16'h0);
  assign T4224 = T4225 ? 5'h1f : 5'h0;
  assign T4225 = T4222[6'h29:6'h29];
  assign twiddle4_3_169_imag = T4228 + T4226;
  assign T4226 = $signed(T4227) / $signed(22'h100000);
  assign T4227 = $signed(31'h3ffe1287) * $signed(16'hffff);
  assign T4228 = {T4231, T4229};
  assign T4229 = $signed(T4230) / $signed(22'h100000);
  assign T4230 = $signed(25'hfb514b) * $signed(16'h0);
  assign T4231 = T4232 ? 6'h3f : 6'h0;
  assign T4232 = T4229[6'h28:6'h28];
  assign T4233 = T2943[1'h0:1'h0];
  assign T4234 = T4249 ? twiddle4_3_171_imag : twiddle4_3_170_imag;
  assign twiddle4_3_170_imag = T4237 + T4235;
  assign T4235 = $signed(T4236) / $signed(22'h100000);
  assign T4236 = $signed(31'h3fffb10b) * $signed(16'hffff);
  assign T4237 = {T4240, T4238};
  assign T4238 = $signed(T4239) / $signed(22'h100000);
  assign T4239 = $signed(24'h6487c3) * $signed(16'h0);
  assign T4240 = T4241 ? 7'h7f : 7'h0;
  assign T4241 = T4238[6'h27:6'h27];
  assign twiddle4_3_171_imag = T4244 + T4242;
  assign T4242 = $signed(T4243) / $signed(22'h100000);
  assign T4243 = $signed(31'h3fffec42) * $signed(16'hffff);
  assign T4244 = {T4247, T4245};
  assign T4245 = $signed(T4246) / $signed(22'h100000);
  assign T4246 = $signed(23'h4dbc0f) * $signed(16'h0);
  assign T4247 = T4248 ? 8'hff : 8'h0;
  assign T4248 = T4245[6'h26:6'h26];
  assign T4249 = T2943[1'h0:1'h0];
  assign T4250 = T2943[1'h1:1'h1];
  assign T4251 = T4284 ? T4268 : T4252;
  assign T4252 = T4267 ? twiddle4_3_173_imag : twiddle4_3_172_imag;
  assign twiddle4_3_172_imag = T4255 + T4253;
  assign T4253 = $signed(T4254) / $signed(22'h100000);
  assign T4254 = $signed(31'h3ffec42d) * $signed(16'hffff);
  assign T4255 = {T4258, T4256};
  assign T4256 = $signed(T4257) / $signed(22'h100000);
  assign T4257 = $signed(25'h136f171) * $signed(16'h0);
  assign T4258 = T4259 ? 6'h3f : 6'h0;
  assign T4259 = T4256[6'h28:6'h28];
  assign twiddle4_3_173_imag = T4262 + T4260;
  assign T4260 = $signed(T4261) / $signed(22'h100000);
  assign T4261 = $signed(31'h3ffc38d0) * $signed(16'hffff);
  assign T4262 = {T4265, T4263};
  assign T4263 = $signed(T4264) / $signed(22'h100000);
  assign T4264 = $signed(26'h2a02b2e) * $signed(16'h0);
  assign T4265 = T4266 ? 5'h1f : 5'h0;
  assign T4266 = T4263[6'h29:6'h29];
  assign T4267 = T2943[1'h0:1'h0];
  assign T4268 = T4283 ? twiddle4_3_175_imag : twiddle4_3_174_imag;
  assign twiddle4_3_174_imag = T4271 + T4269;
  assign T4269 = $signed(T4270) / $signed(22'h100000);
  assign T4270 = $signed(31'h3ff84a3b) * $signed(16'hffff);
  assign T4271 = {T4274, T4272};
  assign T4272 = $signed(T4273) / $signed(22'h100000);
  assign T4273 = $signed(26'h2096c8d) * $signed(16'h0);
  assign T4274 = T4275 ? 5'h1f : 5'h0;
  assign T4275 = T4272[6'h29:6'h29];
  assign twiddle4_3_175_imag = T4278 + T4276;
  assign T4276 = $signed(T4277) / $signed(22'h100000);
  assign T4277 = $signed(31'h3ff2f884) * $signed(16'hffff);
  assign T4278 = {T4281, T4279};
  assign T4279 = $signed(T4280) / $signed(22'h100000);
  assign T4280 = $signed(27'h572b8d3) * $signed(16'h0);
  assign T4281 = T4282 ? 4'hf : 4'h0;
  assign T4282 = T4279[6'h2a:6'h2a];
  assign T4283 = T2943[1'h0:1'h0];
  assign T4284 = T2943[1'h1:1'h1];
  assign T4285 = T2943[2'h2:2'h2];
  assign T4286 = T2943[2'h3:2'h3];
  assign T4287 = T4428 ? T4358 : T4288;
  assign T4288 = T4357 ? T4323 : T4289;
  assign T4289 = T4322 ? T4306 : T4290;
  assign T4290 = T4305 ? twiddle4_3_177_imag : twiddle4_3_176_imag;
  assign twiddle4_3_176_imag = T4293 + T4291;
  assign T4291 = $signed(T4292) / $signed(22'h100000);
  assign T4292 = $signed(31'h3fec43c6) * $signed(16'hffff);
  assign T4293 = {T4296, T4294};
  assign T4294 = $signed(T4295) / $signed(22'h100000);
  assign T4295 = $signed(27'h4dc1342) * $signed(16'h0);
  assign T4296 = T4297 ? 4'hf : 4'h0;
  assign T4297 = T4294[6'h2a:6'h2a];
  assign twiddle4_3_177_imag = T4300 + T4298;
  assign T4298 = $signed(T4299) / $signed(22'h100000);
  assign T4299 = $signed(31'h3fe42c29) * $signed(16'hffff);
  assign T4300 = {T4303, T4301};
  assign T4301 = $signed(T4302) / $signed(22'h100000);
  assign T4302 = $signed(27'h4457f21) * $signed(16'h0);
  assign T4303 = T4304 ? 4'hf : 4'h0;
  assign T4304 = T4301[6'h2a:6'h2a];
  assign T4305 = T2943[1'h0:1'h0];
  assign T4306 = T4321 ? twiddle4_3_179_imag : twiddle4_3_178_imag;
  assign twiddle4_3_178_imag = T4309 + T4307;
  assign T4307 = $signed(T4308) / $signed(22'h100000);
  assign T4308 = $signed(31'h3fdab1d9) * $signed(16'hffff);
  assign T4309 = {T4312, T4310};
  assign T4310 = $signed(T4311) / $signed(22'h100000);
  assign T4311 = $signed(28'hbaeffb3) * $signed(16'h0);
  assign T4312 = T4313 ? 3'h7 : 3'h0;
  assign T4313 = T4310[6'h2b:6'h2b];
  assign twiddle4_3_179_imag = T4316 + T4314;
  assign T4314 = $signed(T4315) / $signed(22'h100000);
  assign T4315 = $signed(31'h3fcfd50a) * $signed(16'hffff);
  assign T4316 = {T4319, T4317};
  assign T4317 = $signed(T4318) / $signed(22'h100000);
  assign T4318 = $signed(28'hb18983c) * $signed(16'h0);
  assign T4319 = T4320 ? 3'h7 : 3'h0;
  assign T4320 = T4317[6'h2b:6'h2b];
  assign T4321 = T2943[1'h0:1'h0];
  assign T4322 = T2943[1'h1:1'h1];
  assign T4323 = T4356 ? T4340 : T4324;
  assign T4324 = T4339 ? twiddle4_3_181_imag : twiddle4_3_180_imag;
  assign twiddle4_3_180_imag = T4327 + T4325;
  assign T4325 = $signed(T4326) / $signed(22'h100000);
  assign T4326 = $signed(31'h3fc395f9) * $signed(16'hffff);
  assign T4327 = {T4330, T4328};
  assign T4328 = $signed(T4329) / $signed(22'h100000);
  assign T4329 = $signed(28'ha824bfe) * $signed(16'h0);
  assign T4330 = T4331 ? 3'h7 : 3'h0;
  assign T4331 = T4328[6'h2b:6'h2b];
  assign twiddle4_3_181_imag = T4334 + T4332;
  assign T4332 = $signed(T4333) / $signed(22'h100000);
  assign T4333 = $signed(31'h3fb5f4ea) * $signed(16'hffff);
  assign T4334 = {T4337, T4335};
  assign T4335 = $signed(T4336) / $signed(22'h100000);
  assign T4336 = $signed(28'h9ec1e3c) * $signed(16'h0);
  assign T4337 = T4338 ? 3'h7 : 3'h0;
  assign T4338 = T4335[6'h2b:6'h2b];
  assign T4339 = T2943[1'h0:1'h0];
  assign T4340 = T4355 ? twiddle4_3_183_imag : twiddle4_3_182_imag;
  assign twiddle4_3_182_imag = T4343 + T4341;
  assign T4341 = $signed(T4342) / $signed(22'h100000);
  assign T4342 = $signed(31'h3fa6f228) * $signed(16'hffff);
  assign T4343 = {T4346, T4344};
  assign T4344 = $signed(T4345) / $signed(22'h100000);
  assign T4345 = $signed(28'h9561237) * $signed(16'h0);
  assign T4346 = T4347 ? 3'h7 : 3'h0;
  assign T4347 = T4344[6'h2b:6'h2b];
  assign twiddle4_3_183_imag = T4350 + T4348;
  assign T4348 = $signed(T4349) / $signed(22'h100000);
  assign T4349 = $signed(31'h3f968e07) * $signed(16'hffff);
  assign T4350 = {T4353, T4351};
  assign T4351 = $signed(T4352) / $signed(22'h100000);
  assign T4352 = $signed(28'h8c02b32) * $signed(16'h0);
  assign T4353 = T4354 ? 3'h7 : 3'h0;
  assign T4354 = T4351[6'h2b:6'h2b];
  assign T4355 = T2943[1'h0:1'h0];
  assign T4356 = T2943[1'h1:1'h1];
  assign T4357 = T2943[2'h2:2'h2];
  assign T4358 = T4427 ? T4393 : T4359;
  assign T4359 = T4392 ? T4376 : T4360;
  assign T4360 = T4375 ? twiddle4_3_185_imag : twiddle4_3_184_imag;
  assign twiddle4_3_184_imag = T4363 + T4361;
  assign T4361 = $signed(T4362) / $signed(22'h100000);
  assign T4362 = $signed(31'h3f84c8e1) * $signed(16'hffff);
  assign T4363 = {T4366, T4364};
  assign T4364 = $signed(T4365) / $signed(22'h100000);
  assign T4365 = $signed(28'h82a6c6b) * $signed(16'h0);
  assign T4366 = T4367 ? 3'h7 : 3'h0;
  assign T4367 = T4364[6'h2b:6'h2b];
  assign twiddle4_3_185_imag = T4370 + T4368;
  assign T4368 = $signed(T4369) / $signed(22'h100000);
  assign T4369 = $signed(31'h3f71a31a) * $signed(16'hffff);
  assign T4370 = {T4373, T4371};
  assign T4371 = $signed(T4372) / $signed(22'h100000);
  assign T4372 = $signed(29'h1794d922) * $signed(16'h0);
  assign T4373 = T4374 ? 2'h3 : 2'h0;
  assign T4374 = T4371[6'h2c:6'h2c];
  assign T4375 = T2943[1'h0:1'h0];
  assign T4376 = T4391 ? twiddle4_3_187_imag : twiddle4_3_186_imag;
  assign twiddle4_3_186_imag = T4379 + T4377;
  assign T4377 = $signed(T4378) / $signed(22'h100000);
  assign T4378 = $signed(31'h3f5d1d1c) * $signed(16'hffff);
  assign T4379 = {T4382, T4380};
  assign T4380 = $signed(T4381) / $signed(22'h100000);
  assign T4381 = $signed(29'h16ff7496) * $signed(16'h0);
  assign T4382 = T4383 ? 2'h3 : 2'h0;
  assign T4383 = T4380[6'h2c:6'h2c];
  assign twiddle4_3_187_imag = T4386 + T4384;
  assign T4384 = $signed(T4385) / $signed(22'h100000);
  assign T4385 = $signed(31'h3f473758) * $signed(16'hffff);
  assign T4386 = {T4389, T4387};
  assign T4387 = $signed(T4388) / $signed(22'h100000);
  assign T4388 = $signed(29'h166a4204) * $signed(16'h0);
  assign T4389 = T4390 ? 2'h3 : 2'h0;
  assign T4390 = T4387[6'h2c:6'h2c];
  assign T4391 = T2943[1'h0:1'h0];
  assign T4392 = T2943[1'h1:1'h1];
  assign T4393 = T4426 ? T4410 : T4394;
  assign T4394 = T4409 ? twiddle4_3_189_imag : twiddle4_3_188_imag;
  assign twiddle4_3_188_imag = T4397 + T4395;
  assign T4395 = $signed(T4396) / $signed(22'h100000);
  assign T4396 = $signed(31'h3f2ff249) * $signed(16'hffff);
  assign T4397 = {T4400, T4398};
  assign T4398 = $signed(T4399) / $signed(22'h100000);
  assign T4399 = $signed(29'h15d544a8) * $signed(16'h0);
  assign T4400 = T4401 ? 2'h3 : 2'h0;
  assign T4401 = T4398[6'h2c:6'h2c];
  assign twiddle4_3_189_imag = T4404 + T4402;
  assign T4402 = $signed(T4403) / $signed(22'h100000);
  assign T4403 = $signed(31'h3f174e6f) * $signed(16'hffff);
  assign T4404 = {T4407, T4405};
  assign T4405 = $signed(T4406) / $signed(22'h100000);
  assign T4406 = $signed(29'h15407fbd) * $signed(16'h0);
  assign T4407 = T4408 ? 2'h3 : 2'h0;
  assign T4408 = T4405[6'h2c:6'h2c];
  assign T4409 = T2943[1'h0:1'h0];
  assign T4410 = T4425 ? twiddle4_3_191_imag : twiddle4_3_190_imag;
  assign twiddle4_3_190_imag = T4413 + T4411;
  assign T4411 = $signed(T4412) / $signed(22'h100000);
  assign T4412 = $signed(31'h3efd4c53) * $signed(16'hffff);
  assign T4413 = {T4416, T4414};
  assign T4414 = $signed(T4415) / $signed(22'h100000);
  assign T4415 = $signed(29'h14abf67e) * $signed(16'h0);
  assign T4416 = T4417 ? 2'h3 : 2'h0;
  assign T4417 = T4414[6'h2c:6'h2c];
  assign twiddle4_3_191_imag = T4420 + T4418;
  assign T4418 = $signed(T4419) / $signed(22'h100000);
  assign T4419 = $signed(31'h3ee1ec86) * $signed(16'hffff);
  assign T4420 = {T4423, T4421};
  assign T4421 = $signed(T4422) / $signed(22'h100000);
  assign T4422 = $signed(29'h1417ac23) * $signed(16'h0);
  assign T4423 = T4424 ? 2'h3 : 2'h0;
  assign T4424 = T4421[6'h2c:6'h2c];
  assign T4425 = T2943[1'h0:1'h0];
  assign T4426 = T2943[1'h1:1'h1];
  assign T4427 = T2943[2'h2:2'h2];
  assign T4428 = T2943[2'h3:2'h3];
  assign T4429 = T2943[3'h4:3'h4];
  assign T4430 = T2943[3'h5:3'h5];
  assign T4431 = T4891 ? T4693 : T4432;
  assign T4432 = T4692 ? T4566 : T4433;
  assign T4433 = T4565 ? T4503 : T4434;
  assign T4434 = T4502 ? T4469 : T4435;
  assign T4435 = T4468 ? T4452 : T4436;
  assign T4436 = T4451 ? twiddle4_3_193_imag : twiddle4_3_192_imag;
  assign twiddle4_3_192_imag = T4439 + T4437;
  assign T4437 = $signed(T4438) / $signed(22'h100000);
  assign T4438 = $signed(31'h3ec52f9f) * $signed(16'hffff);
  assign T4439 = {T4442, T4440};
  assign T4440 = $signed(T4441) / $signed(22'h100000);
  assign T4441 = $signed(29'h1383a3e2) * $signed(16'h0);
  assign T4442 = T4443 ? 2'h3 : 2'h0;
  assign T4443 = T4440[6'h2c:6'h2c];
  assign twiddle4_3_193_imag = T4446 + T4444;
  assign T4444 = $signed(T4445) / $signed(22'h100000);
  assign T4445 = $signed(31'h3ea7163f) * $signed(16'hffff);
  assign T4446 = {T4449, T4447};
  assign T4447 = $signed(T4448) / $signed(22'h100000);
  assign T4448 = $signed(29'h12efe0f3) * $signed(16'h0);
  assign T4449 = T4450 ? 2'h3 : 2'h0;
  assign T4450 = T4447[6'h2c:6'h2c];
  assign T4451 = T2943[1'h0:1'h0];
  assign T4452 = T4467 ? twiddle4_3_195_imag : twiddle4_3_194_imag;
  assign twiddle4_3_194_imag = T4455 + T4453;
  assign T4453 = $signed(T4454) / $signed(22'h100000);
  assign T4454 = $signed(31'h3e87a10b) * $signed(16'hffff);
  assign T4455 = {T4458, T4456};
  assign T4456 = $signed(T4457) / $signed(22'h100000);
  assign T4457 = $signed(29'h125c6689) * $signed(16'h0);
  assign T4458 = T4459 ? 2'h3 : 2'h0;
  assign T4459 = T4456[6'h2c:6'h2c];
  assign twiddle4_3_195_imag = T4462 + T4460;
  assign T4460 = $signed(T4461) / $signed(22'h100000);
  assign T4461 = $signed(31'h3e66d0b4) * $signed(16'hffff);
  assign T4462 = {T4465, T4463};
  assign T4463 = $signed(T4464) / $signed(22'h100000);
  assign T4464 = $signed(29'h11c937d7) * $signed(16'h0);
  assign T4465 = T4466 ? 2'h3 : 2'h0;
  assign T4466 = T4463[6'h2c:6'h2c];
  assign T4467 = T2943[1'h0:1'h0];
  assign T4468 = T2943[1'h1:1'h1];
  assign T4469 = T4501 ? T4486 : T4470;
  assign T4470 = T4485 ? twiddle4_3_197_imag : twiddle4_3_196_imag;
  assign twiddle4_3_196_imag = T4473 + T4471;
  assign T4471 = $signed(T4472) / $signed(22'h100000);
  assign T4472 = $signed(31'h3e44a5ee) * $signed(16'hffff);
  assign T4473 = {T4476, T4474};
  assign T4474 = $signed(T4475) / $signed(22'h100000);
  assign T4475 = $signed(29'h1136580e) * $signed(16'h0);
  assign T4476 = T4477 ? 2'h3 : 2'h0;
  assign T4477 = T4474[6'h2c:6'h2c];
  assign twiddle4_3_197_imag = T4480 + T4478;
  assign T4478 = $signed(T4479) / $signed(22'h100000);
  assign T4479 = $signed(31'h3e212179) * $signed(16'hffff);
  assign T4480 = {T4483, T4481};
  assign T4481 = $signed(T4482) / $signed(22'h100000);
  assign T4482 = $signed(29'h10a3ca5d) * $signed(16'h0);
  assign T4483 = T4484 ? 2'h3 : 2'h0;
  assign T4484 = T4481[6'h2c:6'h2c];
  assign T4485 = T2943[1'h0:1'h0];
  assign T4486 = T4500 ? twiddle4_3_199_imag : twiddle4_3_198_imag;
  assign twiddle4_3_198_imag = T4489 + T4487;
  assign T4487 = $signed(T4488) / $signed(22'h100000);
  assign T4488 = $signed(31'h3dfc4418) * $signed(16'hffff);
  assign T4489 = {T4492, T4490};
  assign T4490 = $signed(T4491) / $signed(22'h100000);
  assign T4491 = $signed(29'h101191f3) * $signed(16'h0);
  assign T4492 = T4493 ? 2'h3 : 2'h0;
  assign T4493 = T4490[6'h2c:6'h2c];
  assign twiddle4_3_199_imag = T4496 + T4494;
  assign T4494 = $signed(T4495) / $signed(22'h100000);
  assign T4495 = $signed(31'h3dd60e98) * $signed(16'hffff);
  assign T4496 = {T4499, T4497};
  assign T4497 = $signed(T4498) / $signed(22'h100000);
  assign T4498 = $signed(30'h2f7fb1fb) * $signed(16'h0);
  assign T4499 = T4497[6'h2d:6'h2d];
  assign T4500 = T2943[1'h0:1'h0];
  assign T4501 = T2943[1'h1:1'h1];
  assign T4502 = T2943[2'h2:2'h2];
  assign T4503 = T4564 ? T4534 : T4504;
  assign T4504 = T4533 ? T4519 : T4505;
  assign T4505 = T4518 ? twiddle4_3_201_imag : twiddle4_3_200_imag;
  assign twiddle4_3_200_imag = T4508 + T4506;
  assign T4506 = $signed(T4507) / $signed(22'h100000);
  assign T4507 = $signed(31'h3dae81ce) * $signed(16'hffff);
  assign T4508 = {T4511, T4509};
  assign T4509 = $signed(T4510) / $signed(22'h100000);
  assign T4510 = $signed(30'h2eee2d9e) * $signed(16'h0);
  assign T4511 = T4509[6'h2d:6'h2d];
  assign twiddle4_3_201_imag = T4514 + T4512;
  assign T4512 = $signed(T4513) / $signed(22'h100000);
  assign T4513 = $signed(31'h3d859e96) * $signed(16'hffff);
  assign T4514 = {T4517, T4515};
  assign T4515 = $signed(T4516) / $signed(22'h100000);
  assign T4516 = $signed(30'h2e5d0805) * $signed(16'h0);
  assign T4517 = T4515[6'h2d:6'h2d];
  assign T4518 = T2943[1'h0:1'h0];
  assign T4519 = T4532 ? twiddle4_3_203_imag : twiddle4_3_202_imag;
  assign twiddle4_3_202_imag = T4522 + T4520;
  assign T4520 = $signed(T4521) / $signed(22'h100000);
  assign T4521 = $signed(31'h3d5b65d1) * $signed(16'hffff);
  assign T4522 = {T4525, T4523};
  assign T4523 = $signed(T4524) / $signed(22'h100000);
  assign T4524 = $signed(30'h2dcc4455) * $signed(16'h0);
  assign T4525 = T4523[6'h2d:6'h2d];
  assign twiddle4_3_203_imag = T4528 + T4526;
  assign T4526 = $signed(T4527) / $signed(22'h100000);
  assign T4527 = $signed(31'h3d2fd86c) * $signed(16'hffff);
  assign T4528 = {T4531, T4529};
  assign T4529 = $signed(T4530) / $signed(22'h100000);
  assign T4530 = $signed(30'h2d3be5b2) * $signed(16'h0);
  assign T4531 = T4529[6'h2d:6'h2d];
  assign T4532 = T2943[1'h0:1'h0];
  assign T4533 = T2943[1'h1:1'h1];
  assign T4534 = T4563 ? T4549 : T4535;
  assign T4535 = T4548 ? twiddle4_3_205_imag : twiddle4_3_204_imag;
  assign twiddle4_3_204_imag = T4538 + T4536;
  assign T4536 = $signed(T4537) / $signed(22'h100000);
  assign T4537 = $signed(31'h3d02f756) * $signed(16'hffff);
  assign T4538 = {T4541, T4539};
  assign T4539 = $signed(T4540) / $signed(22'h100000);
  assign T4540 = $signed(30'h2cabef3e) * $signed(16'h0);
  assign T4541 = T4539[6'h2d:6'h2d];
  assign twiddle4_3_205_imag = T4544 + T4542;
  assign T4542 = $signed(T4543) / $signed(22'h100000);
  assign T4543 = $signed(31'h3cd4c38a) * $signed(16'hffff);
  assign T4544 = {T4547, T4545};
  assign T4545 = $signed(T4546) / $signed(22'h100000);
  assign T4546 = $signed(30'h2c1c6417) * $signed(16'h0);
  assign T4547 = T4545[6'h2d:6'h2d];
  assign T4548 = T2943[1'h0:1'h0];
  assign T4549 = T4562 ? twiddle4_3_207_imag : twiddle4_3_206_imag;
  assign twiddle4_3_206_imag = T4552 + T4550;
  assign T4550 = $signed(T4551) / $signed(22'h100000);
  assign T4551 = $signed(31'h3ca53e08) * $signed(16'hffff);
  assign T4552 = {T4555, T4553};
  assign T4553 = $signed(T4554) / $signed(22'h100000);
  assign T4554 = $signed(30'h2b8d475b) * $signed(16'h0);
  assign T4555 = T4553[6'h2d:6'h2d];
  assign twiddle4_3_207_imag = T4558 + T4556;
  assign T4556 = $signed(T4557) / $signed(22'h100000);
  assign T4557 = $signed(31'h3c7467d8) * $signed(16'hffff);
  assign T4558 = {T4561, T4559};
  assign T4559 = $signed(T4560) / $signed(22'h100000);
  assign T4560 = $signed(30'h2afe9c24) * $signed(16'h0);
  assign T4561 = T4559[6'h2d:6'h2d];
  assign T4562 = T2943[1'h0:1'h0];
  assign T4563 = T2943[1'h1:1'h1];
  assign T4564 = T2943[2'h2:2'h2];
  assign T4565 = T2943[2'h3:2'h3];
  assign T4566 = T4691 ? T4629 : T4567;
  assign T4567 = T4628 ? T4598 : T4568;
  assign T4568 = T4597 ? T4583 : T4569;
  assign T4569 = T4582 ? twiddle4_3_209_imag : twiddle4_3_208_imag;
  assign twiddle4_3_208_imag = T4572 + T4570;
  assign T4570 = $signed(T4571) / $signed(22'h100000);
  assign T4571 = $signed(31'h3c424209) * $signed(16'hffff);
  assign T4572 = {T4575, T4573};
  assign T4573 = $signed(T4574) / $signed(22'h100000);
  assign T4574 = $signed(30'h2a70658b) * $signed(16'h0);
  assign T4575 = T4573[6'h2d:6'h2d];
  assign twiddle4_3_209_imag = T4578 + T4576;
  assign T4576 = $signed(T4577) / $signed(22'h100000);
  assign T4577 = $signed(31'h3c0ecdb2) * $signed(16'hffff);
  assign T4578 = {T4581, T4579};
  assign T4579 = $signed(T4580) / $signed(22'h100000);
  assign T4580 = $signed(30'h29e2a6a4) * $signed(16'h0);
  assign T4581 = T4579[6'h2d:6'h2d];
  assign T4582 = T2943[1'h0:1'h0];
  assign T4583 = T4596 ? twiddle4_3_211_imag : twiddle4_3_210_imag;
  assign twiddle4_3_210_imag = T4586 + T4584;
  assign T4584 = $signed(T4585) / $signed(22'h100000);
  assign T4585 = $signed(31'h3bda0bef) * $signed(16'hffff);
  assign T4586 = {T4589, T4587};
  assign T4587 = $signed(T4588) / $signed(22'h100000);
  assign T4588 = $signed(30'h29556283) * $signed(16'h0);
  assign T4589 = T4587[6'h2d:6'h2d];
  assign twiddle4_3_211_imag = T4592 + T4590;
  assign T4590 = $signed(T4591) / $signed(22'h100000);
  assign T4591 = $signed(31'h3ba3fde7) * $signed(16'hffff);
  assign T4592 = {T4595, T4593};
  assign T4593 = $signed(T4594) / $signed(22'h100000);
  assign T4594 = $signed(30'h28c89c37) * $signed(16'h0);
  assign T4595 = T4593[6'h2d:6'h2d];
  assign T4596 = T2943[1'h0:1'h0];
  assign T4597 = T2943[1'h1:1'h1];
  assign T4598 = T4627 ? T4613 : T4599;
  assign T4599 = T4612 ? twiddle4_3_213_imag : twiddle4_3_212_imag;
  assign twiddle4_3_212_imag = T4602 + T4600;
  assign T4600 = $signed(T4601) / $signed(22'h100000);
  assign T4601 = $signed(31'h3b6ca4c4) * $signed(16'hffff);
  assign T4602 = {T4605, T4603};
  assign T4603 = $signed(T4604) / $signed(22'h100000);
  assign T4604 = $signed(30'h283c56cf) * $signed(16'h0);
  assign T4605 = T4603[6'h2d:6'h2d];
  assign twiddle4_3_213_imag = T4608 + T4606;
  assign T4606 = $signed(T4607) / $signed(22'h100000);
  assign T4607 = $signed(31'h3b3401bb) * $signed(16'hffff);
  assign T4608 = {T4611, T4609};
  assign T4609 = $signed(T4610) / $signed(22'h100000);
  assign T4610 = $signed(30'h27b09556) * $signed(16'h0);
  assign T4611 = T4609[6'h2d:6'h2d];
  assign T4612 = T2943[1'h0:1'h0];
  assign T4613 = T4626 ? twiddle4_3_215_imag : twiddle4_3_214_imag;
  assign twiddle4_3_214_imag = T4616 + T4614;
  assign T4614 = $signed(T4615) / $signed(22'h100000);
  assign T4615 = $signed(31'h3afa1605) * $signed(16'hffff);
  assign T4616 = {T4619, T4617};
  assign T4617 = $signed(T4618) / $signed(22'h100000);
  assign T4618 = $signed(30'h27255ad2) * $signed(16'h0);
  assign T4619 = T4617[6'h2d:6'h2d];
  assign twiddle4_3_215_imag = T4622 + T4620;
  assign T4620 = $signed(T4621) / $signed(22'h100000);
  assign T4621 = $signed(31'h3abee2e5) * $signed(16'hffff);
  assign T4622 = {T4625, T4623};
  assign T4623 = $signed(T4624) / $signed(22'h100000);
  assign T4624 = $signed(30'h269aaa49) * $signed(16'h0);
  assign T4625 = T4623[6'h2d:6'h2d];
  assign T4626 = T2943[1'h0:1'h0];
  assign T4627 = T2943[1'h1:1'h1];
  assign T4628 = T2943[2'h2:2'h2];
  assign T4629 = T4690 ? T4660 : T4630;
  assign T4630 = T4659 ? T4645 : T4631;
  assign T4631 = T4644 ? twiddle4_3_217_imag : twiddle4_3_216_imag;
  assign twiddle4_3_216_imag = T4634 + T4632;
  assign T4632 = $signed(T4633) / $signed(22'h100000);
  assign T4633 = $signed(31'h3a8269a2) * $signed(16'hffff);
  assign T4634 = {T4637, T4635};
  assign T4635 = $signed(T4636) / $signed(22'h100000);
  assign T4636 = $signed(30'h261086bd) * $signed(16'h0);
  assign T4637 = T4635[6'h2d:6'h2d];
  assign twiddle4_3_217_imag = T4640 + T4638;
  assign T4638 = $signed(T4639) / $signed(22'h100000);
  assign T4639 = $signed(31'h3a44ab8d) * $signed(16'hffff);
  assign T4640 = {T4643, T4641};
  assign T4641 = $signed(T4642) / $signed(22'h100000);
  assign T4642 = $signed(30'h2586f32d) * $signed(16'h0);
  assign T4643 = T4641[6'h2d:6'h2d];
  assign T4644 = T2943[1'h0:1'h0];
  assign T4645 = T4658 ? twiddle4_3_219_imag : twiddle4_3_218_imag;
  assign twiddle4_3_218_imag = T4648 + T4646;
  assign T4646 = $signed(T4647) / $signed(22'h100000);
  assign T4647 = $signed(31'h3a05a9fd) * $signed(16'hffff);
  assign T4648 = {T4651, T4649};
  assign T4649 = $signed(T4650) / $signed(22'h100000);
  assign T4650 = $signed(30'h24fdf294) * $signed(16'h0);
  assign T4651 = T4649[6'h2d:6'h2d];
  assign twiddle4_3_219_imag = T4654 + T4652;
  assign T4652 = $signed(T4653) / $signed(22'h100000);
  assign T4653 = $signed(31'h39c5664f) * $signed(16'hffff);
  assign T4654 = {T4657, T4655};
  assign T4655 = $signed(T4656) / $signed(22'h100000);
  assign T4656 = $signed(30'h247587ec) * $signed(16'h0);
  assign T4657 = T4655[6'h2d:6'h2d];
  assign T4658 = T2943[1'h0:1'h0];
  assign T4659 = T2943[1'h1:1'h1];
  assign T4660 = T4689 ? T4675 : T4661;
  assign T4661 = T4674 ? twiddle4_3_221_imag : twiddle4_3_220_imag;
  assign twiddle4_3_220_imag = T4664 + T4662;
  assign T4662 = $signed(T4663) / $signed(22'h100000);
  assign T4663 = $signed(31'h3983e1e7) * $signed(16'hffff);
  assign T4664 = {T4667, T4665};
  assign T4665 = $signed(T4666) / $signed(22'h100000);
  assign T4666 = $signed(30'h23edb628) * $signed(16'h0);
  assign T4667 = T4665[6'h2d:6'h2d];
  assign twiddle4_3_221_imag = T4670 + T4668;
  assign T4668 = $signed(T4669) / $signed(22'h100000);
  assign T4669 = $signed(31'h39411e33) * $signed(16'hffff);
  assign T4670 = {T4673, T4671};
  assign T4671 = $signed(T4672) / $signed(22'h100000);
  assign T4672 = $signed(30'h2366803d) * $signed(16'h0);
  assign T4673 = T4671[6'h2d:6'h2d];
  assign T4674 = T2943[1'h0:1'h0];
  assign T4675 = T4688 ? twiddle4_3_223_imag : twiddle4_3_222_imag;
  assign twiddle4_3_222_imag = T4678 + T4676;
  assign T4676 = $signed(T4677) / $signed(22'h100000);
  assign T4677 = $signed(31'h38fd1ca4) * $signed(16'hffff);
  assign T4678 = {T4681, T4679};
  assign T4679 = $signed(T4680) / $signed(22'h100000);
  assign T4680 = $signed(30'h22dfe918) * $signed(16'h0);
  assign T4681 = T4679[6'h2d:6'h2d];
  assign twiddle4_3_223_imag = T4684 + T4682;
  assign T4682 = $signed(T4683) / $signed(22'h100000);
  assign T4683 = $signed(31'h38b7deb3) * $signed(16'hffff);
  assign T4684 = {T4687, T4685};
  assign T4685 = $signed(T4686) / $signed(22'h100000);
  assign T4686 = $signed(30'h2259f3a4) * $signed(16'h0);
  assign T4687 = T4685[6'h2d:6'h2d];
  assign T4688 = T2943[1'h0:1'h0];
  assign T4689 = T2943[1'h1:1'h1];
  assign T4690 = T2943[2'h2:2'h2];
  assign T4691 = T2943[2'h3:2'h3];
  assign T4692 = T2943[3'h4:3'h4];
  assign T4693 = T4890 ? T4796 : T4694;
  assign T4694 = T4795 ? T4749 : T4695;
  assign T4695 = T4748 ? T4726 : T4696;
  assign T4696 = T4725 ? T4711 : T4697;
  assign T4697 = T4710 ? twiddle4_3_225_imag : twiddle4_3_224_imag;
  assign twiddle4_3_224_imag = T4700 + T4698;
  assign T4698 = $signed(T4699) / $signed(22'h100000);
  assign T4699 = $signed(31'h387165e3) * $signed(16'hffff);
  assign T4700 = {T4703, T4701};
  assign T4701 = $signed(T4702) / $signed(22'h100000);
  assign T4702 = $signed(30'h21d4a2c8) * $signed(16'h0);
  assign T4703 = T4701[6'h2d:6'h2d];
  assign twiddle4_3_225_imag = T4706 + T4704;
  assign T4704 = $signed(T4705) / $signed(22'h100000);
  assign T4705 = $signed(31'h3829b3b8) * $signed(16'hffff);
  assign T4706 = {T4709, T4707};
  assign T4707 = $signed(T4708) / $signed(22'h100000);
  assign T4708 = $signed(30'h214ff96b) * $signed(16'h0);
  assign T4709 = T4707[6'h2d:6'h2d];
  assign T4710 = T2943[1'h0:1'h0];
  assign T4711 = T4724 ? twiddle4_3_227_imag : twiddle4_3_226_imag;
  assign twiddle4_3_226_imag = T4714 + T4712;
  assign T4712 = $signed(T4713) / $signed(22'h100000);
  assign T4713 = $signed(31'h37e0c9c2) * $signed(16'hffff);
  assign T4714 = {T4717, T4715};
  assign T4715 = $signed(T4716) / $signed(22'h100000);
  assign T4716 = $signed(30'h20cbfa6a) * $signed(16'h0);
  assign T4717 = T4715[6'h2d:6'h2d];
  assign twiddle4_3_227_imag = T4720 + T4718;
  assign T4718 = $signed(T4719) / $signed(22'h100000);
  assign T4719 = $signed(31'h3796a996) * $signed(16'hffff);
  assign T4720 = {T4723, T4721};
  assign T4721 = $signed(T4722) / $signed(22'h100000);
  assign T4722 = $signed(30'h2048a8a4) * $signed(16'h0);
  assign T4723 = T4721[6'h2d:6'h2d];
  assign T4724 = T2943[1'h0:1'h0];
  assign T4725 = T2943[1'h1:1'h1];
  assign T4726 = T4747 ? T4737 : T4727;
  assign T4727 = T4736 ? twiddle4_3_229_imag : twiddle4_3_228_imag;
  assign twiddle4_3_228_imag = T4730 + T4728;
  assign T4728 = $signed(T4729) / $signed(22'h100000);
  assign T4729 = $signed(31'h374b54ce) * $signed(16'hffff);
  assign T4730 = $signed(T4731) / $signed(22'h100000);
  assign T4731 = $signed(31'h5fc606f2) * $signed(16'h0);
  assign twiddle4_3_229_imag = T4734 + T4732;
  assign T4732 = $signed(T4733) / $signed(22'h100000);
  assign T4733 = $signed(31'h36fecd0d) * $signed(16'hffff);
  assign T4734 = $signed(T4735) / $signed(22'h100000);
  assign T4735 = $signed(31'h5f441828) * $signed(16'h0);
  assign T4736 = T2943[1'h0:1'h0];
  assign T4737 = T4746 ? twiddle4_3_231_imag : twiddle4_3_230_imag;
  assign twiddle4_3_230_imag = T4740 + T4738;
  assign T4738 = $signed(T4739) / $signed(22'h100000);
  assign T4739 = $signed(31'h36b113fd) * $signed(16'hffff);
  assign T4740 = $signed(T4741) / $signed(22'h100000);
  assign T4741 = $signed(31'h5ec2df18) * $signed(16'h0);
  assign twiddle4_3_231_imag = T4744 + T4742;
  assign T4742 = $signed(T4743) / $signed(22'h100000);
  assign T4743 = $signed(31'h36622b4b) * $signed(16'hffff);
  assign T4744 = $signed(T4745) / $signed(22'h100000);
  assign T4745 = $signed(31'h5e425e90) * $signed(16'h0);
  assign T4746 = T2943[1'h0:1'h0];
  assign T4747 = T2943[1'h1:1'h1];
  assign T4748 = T2943[2'h2:2'h2];
  assign T4749 = T4794 ? T4772 : T4750;
  assign T4750 = T4771 ? T4761 : T4751;
  assign T4751 = T4760 ? twiddle4_3_233_imag : twiddle4_3_232_imag;
  assign twiddle4_3_232_imag = T4754 + T4752;
  assign T4752 = $signed(T4753) / $signed(22'h100000);
  assign T4753 = $signed(31'h361214b0) * $signed(16'hffff);
  assign T4754 = $signed(T4755) / $signed(22'h100000);
  assign T4755 = $signed(31'h5dc29958) * $signed(16'h0);
  assign twiddle4_3_233_imag = T4758 + T4756;
  assign T4756 = $signed(T4757) / $signed(22'h100000);
  assign T4757 = $signed(31'h35c0d1e6) * $signed(16'hffff);
  assign T4758 = $signed(T4759) / $signed(22'h100000);
  assign T4759 = $signed(31'h5d439237) * $signed(16'h0);
  assign T4760 = T2943[1'h0:1'h0];
  assign T4761 = T4770 ? twiddle4_3_235_imag : twiddle4_3_234_imag;
  assign twiddle4_3_234_imag = T4764 + T4762;
  assign T4762 = $signed(T4763) / $signed(22'h100000);
  assign T4763 = $signed(31'h356e64b2) * $signed(16'hffff);
  assign T4764 = $signed(T4765) / $signed(22'h100000);
  assign T4765 = $signed(31'h5cc54bed) * $signed(16'h0);
  assign twiddle4_3_235_imag = T4768 + T4766;
  assign T4766 = $signed(T4767) / $signed(22'h100000);
  assign T4767 = $signed(31'h351acedc) * $signed(16'hffff);
  assign T4768 = $signed(T4769) / $signed(22'h100000);
  assign T4769 = $signed(31'h5c47c937) * $signed(16'h0);
  assign T4770 = T2943[1'h0:1'h0];
  assign T4771 = T2943[1'h1:1'h1];
  assign T4772 = T4793 ? T4783 : T4773;
  assign T4773 = T4782 ? twiddle4_3_237_imag : twiddle4_3_236_imag;
  assign twiddle4_3_236_imag = T4776 + T4774;
  assign T4774 = $signed(T4775) / $signed(22'h100000);
  assign T4775 = $signed(31'h34c61236) * $signed(16'hffff);
  assign T4776 = $signed(T4777) / $signed(22'h100000);
  assign T4777 = $signed(31'h5bcb0cce) * $signed(16'h0);
  assign twiddle4_3_237_imag = T4780 + T4778;
  assign T4778 = $signed(T4779) / $signed(22'h100000);
  assign T4779 = $signed(31'h34703094) * $signed(16'hffff);
  assign T4780 = $signed(T4781) / $signed(22'h100000);
  assign T4781 = $signed(31'h5b4f1967) * $signed(16'h0);
  assign T4782 = T2943[1'h0:1'h0];
  assign T4783 = T4792 ? twiddle4_3_239_imag : twiddle4_3_238_imag;
  assign twiddle4_3_238_imag = T4786 + T4784;
  assign T4784 = $signed(T4785) / $signed(22'h100000);
  assign T4785 = $signed(31'h34192bd5) * $signed(16'hffff);
  assign T4786 = $signed(T4787) / $signed(22'h100000);
  assign T4787 = $signed(31'h5ad3f1b2) * $signed(16'h0);
  assign twiddle4_3_239_imag = T4790 + T4788;
  assign T4788 = $signed(T4789) / $signed(22'h100000);
  assign T4789 = $signed(31'h33c105db) * $signed(16'hffff);
  assign T4790 = $signed(T4791) / $signed(22'h100000);
  assign T4791 = $signed(31'h5a59985a) * $signed(16'h0);
  assign T4792 = T2943[1'h0:1'h0];
  assign T4793 = T2943[1'h1:1'h1];
  assign T4794 = T2943[2'h2:2'h2];
  assign T4795 = T2943[2'h3:2'h3];
  assign T4796 = T4889 ? T4843 : T4797;
  assign T4797 = T4842 ? T4820 : T4798;
  assign T4798 = T4819 ? T4809 : T4799;
  assign T4799 = T4808 ? twiddle4_3_241_imag : twiddle4_3_240_imag;
  assign twiddle4_3_240_imag = T4802 + T4800;
  assign T4800 = $signed(T4801) / $signed(22'h100000);
  assign T4801 = $signed(31'h3367c08f) * $signed(16'hffff);
  assign T4802 = $signed(T4803) / $signed(22'h100000);
  assign T4803 = $signed(31'h59e01007) * $signed(16'h0);
  assign twiddle4_3_241_imag = T4806 + T4804;
  assign T4804 = $signed(T4805) / $signed(22'h100000);
  assign T4805 = $signed(31'h330d5de2) * $signed(16'hffff);
  assign T4806 = $signed(T4807) / $signed(22'h100000);
  assign T4807 = $signed(31'h59675b5b) * $signed(16'h0);
  assign T4808 = T2943[1'h0:1'h0];
  assign T4809 = T4818 ? twiddle4_3_243_imag : twiddle4_3_242_imag;
  assign twiddle4_3_242_imag = T4812 + T4810;
  assign T4810 = $signed(T4811) / $signed(22'h100000);
  assign T4811 = $signed(31'h32b1dfc9) * $signed(16'hffff);
  assign T4812 = $signed(T4813) / $signed(22'h100000);
  assign T4813 = $signed(31'h58ef7cf5) * $signed(16'h0);
  assign twiddle4_3_243_imag = T4816 + T4814;
  assign T4814 = $signed(T4815) / $signed(22'h100000);
  assign T4815 = $signed(31'h3255483f) * $signed(16'hffff);
  assign T4816 = $signed(T4817) / $signed(22'h100000);
  assign T4817 = $signed(31'h5878776d) * $signed(16'h0);
  assign T4818 = T2943[1'h0:1'h0];
  assign T4819 = T2943[1'h1:1'h1];
  assign T4820 = T4841 ? T4831 : T4821;
  assign T4821 = T4830 ? twiddle4_3_245_imag : twiddle4_3_244_imag;
  assign twiddle4_3_244_imag = T4824 + T4822;
  assign T4822 = $signed(T4823) / $signed(22'h100000);
  assign T4823 = $signed(31'h31f79947) * $signed(16'hffff);
  assign T4824 = $signed(T4825) / $signed(22'h100000);
  assign T4825 = $signed(31'h58024d5a) * $signed(16'h0);
  assign twiddle4_3_245_imag = T4828 + T4826;
  assign T4826 = $signed(T4827) / $signed(22'h100000);
  assign T4827 = $signed(31'h3198d4ea) * $signed(16'hffff);
  assign T4828 = $signed(T4829) / $signed(22'h100000);
  assign T4829 = $signed(31'h578d014a) * $signed(16'h0);
  assign T4830 = T2943[1'h0:1'h0];
  assign T4831 = T4840 ? twiddle4_3_247_imag : twiddle4_3_246_imag;
  assign twiddle4_3_246_imag = T4834 + T4832;
  assign T4832 = $signed(T4833) / $signed(22'h100000);
  assign T4833 = $signed(31'h3138fd34) * $signed(16'hffff);
  assign T4834 = $signed(T4835) / $signed(22'h100000);
  assign T4835 = $signed(31'h571895c9) * $signed(16'h0);
  assign twiddle4_3_247_imag = T4838 + T4836;
  assign T4836 = $signed(T4837) / $signed(22'h100000);
  assign T4837 = $signed(31'h30d8143b) * $signed(16'hffff);
  assign T4838 = $signed(T4839) / $signed(22'h100000);
  assign T4839 = $signed(31'h56a50d5e) * $signed(16'h0);
  assign T4840 = T2943[1'h0:1'h0];
  assign T4841 = T2943[1'h1:1'h1];
  assign T4842 = T2943[2'h2:2'h2];
  assign T4843 = T4888 ? T4866 : T4844;
  assign T4844 = T4865 ? T4855 : T4845;
  assign T4845 = T4854 ? twiddle4_3_249_imag : twiddle4_3_248_imag;
  assign twiddle4_3_248_imag = T4848 + T4846;
  assign T4846 = $signed(T4847) / $signed(22'h100000);
  assign T4847 = $signed(31'h30761c17) * $signed(16'hffff);
  assign T4848 = $signed(T4849) / $signed(22'h100000);
  assign T4849 = $signed(31'h56326a89) * $signed(16'h0);
  assign twiddle4_3_249_imag = T4852 + T4850;
  assign T4850 = $signed(T4851) / $signed(22'h100000);
  assign T4851 = $signed(31'h301316ea) * $signed(16'hffff);
  assign T4852 = $signed(T4853) / $signed(22'h100000);
  assign T4853 = $signed(31'h55c0afc7) * $signed(16'h0);
  assign T4854 = T2943[1'h0:1'h0];
  assign T4855 = T4864 ? twiddle4_3_251_imag : twiddle4_3_250_imag;
  assign twiddle4_3_250_imag = T4858 + T4856;
  assign T4856 = $signed(T4857) / $signed(22'h100000);
  assign T4857 = $signed(31'h2faf06d9) * $signed(16'hffff);
  assign T4858 = $signed(T4859) / $signed(22'h100000);
  assign T4859 = $signed(31'h554fdf8f) * $signed(16'h0);
  assign twiddle4_3_251_imag = T4862 + T4860;
  assign T4860 = $signed(T4861) / $signed(22'h100000);
  assign T4861 = $signed(31'h2f49ee0f) * $signed(16'hffff);
  assign T4862 = $signed(T4863) / $signed(22'h100000);
  assign T4863 = $signed(31'h54dffc55) * $signed(16'h0);
  assign T4864 = T2943[1'h0:1'h0];
  assign T4865 = T2943[1'h1:1'h1];
  assign T4866 = T4887 ? T4877 : T4867;
  assign T4867 = T4876 ? twiddle4_3_253_imag : twiddle4_3_252_imag;
  assign twiddle4_3_252_imag = T4870 + T4868;
  assign T4868 = $signed(T4869) / $signed(22'h100000);
  assign T4869 = $signed(31'h2ee3cebe) * $signed(16'hffff);
  assign T4870 = $signed(T4871) / $signed(22'h100000);
  assign T4871 = $signed(31'h54710884) * $signed(16'h0);
  assign twiddle4_3_253_imag = T4874 + T4872;
  assign T4872 = $signed(T4873) / $signed(22'h100000);
  assign T4873 = $signed(31'h2e7cab1c) * $signed(16'hffff);
  assign T4874 = $signed(T4875) / $signed(22'h100000);
  assign T4875 = $signed(31'h54030685) * $signed(16'h0);
  assign T4876 = T2943[1'h0:1'h0];
  assign T4877 = T4886 ? twiddle4_3_255_imag : twiddle4_3_254_imag;
  assign twiddle4_3_254_imag = T4880 + T4878;
  assign T4878 = $signed(T4879) / $signed(22'h100000);
  assign T4879 = $signed(31'h2e148566) * $signed(16'hffff);
  assign T4880 = $signed(T4881) / $signed(22'h100000);
  assign T4881 = $signed(31'h5395f8ba) * $signed(16'h0);
  assign twiddle4_3_255_imag = T4884 + T4882;
  assign T4882 = $signed(T4883) / $signed(22'h100000);
  assign T4883 = $signed(31'h2dab5fde) * $signed(16'hffff);
  assign T4884 = $signed(T4885) / $signed(22'h100000);
  assign T4885 = $signed(31'h5329e182) * $signed(16'h0);
  assign T4886 = T2943[1'h0:1'h0];
  assign T4887 = T2943[1'h1:1'h1];
  assign T4888 = T2943[2'h2:2'h2];
  assign T4889 = T2943[2'h3:2'h3];
  assign T4890 = T2943[3'h4:3'h4];
  assign T4891 = T2943[3'h5:3'h5];
  assign T4892 = T2943[3'h6:3'h6];
  assign T4893 = T3872[6'h2e:6'h2e];
  assign T4894 = T2943[3'h7:3'h7];
  assign T4895 = {T6852, T4896};
  assign T4896 = T6851 ? T5916 : T4897;
  assign T4897 = T5915 ? T5356 : T4898;
  assign T4898 = T5355 ? T5095 : T4899;
  assign T4899 = T5094 ? T4994 : T4900;
  assign T4900 = T4993 ? T4947 : T4901;
  assign T4901 = T4946 ? T4924 : T4902;
  assign T4902 = T4923 ? T4913 : T4903;
  assign T4903 = T4912 ? twiddle4_3_257_imag : twiddle4_3_256_imag;
  assign twiddle4_3_256_imag = T4906 + T4904;
  assign T4904 = $signed(T4905) / $signed(22'h100000);
  assign T4905 = $signed(31'h2d413ccc) * $signed(16'hffff);
  assign T4906 = $signed(T4907) / $signed(22'h100000);
  assign T4907 = $signed(31'h52bec334) * $signed(16'h0);
  assign twiddle4_3_257_imag = T4910 + T4908;
  assign T4908 = $signed(T4909) / $signed(22'h100000);
  assign T4909 = $signed(31'h2cd61e7e) * $signed(16'hffff);
  assign T4910 = $signed(T4911) / $signed(22'h100000);
  assign T4911 = $signed(31'h5254a022) * $signed(16'h0);
  assign T4912 = T2943[1'h0:1'h0];
  assign T4913 = T4922 ? twiddle4_3_259_imag : twiddle4_3_258_imag;
  assign twiddle4_3_258_imag = T4916 + T4914;
  assign T4914 = $signed(T4915) / $signed(22'h100000);
  assign T4915 = $signed(31'h2c6a0746) * $signed(16'hffff);
  assign T4916 = $signed(T4917) / $signed(22'h100000);
  assign T4917 = $signed(31'h51eb7a9a) * $signed(16'h0);
  assign twiddle4_3_259_imag = T4920 + T4918;
  assign T4918 = $signed(T4919) / $signed(22'h100000);
  assign T4919 = $signed(31'h2bfcf97b) * $signed(16'hffff);
  assign T4920 = $signed(T4921) / $signed(22'h100000);
  assign T4921 = $signed(31'h518354e4) * $signed(16'h0);
  assign T4922 = T2943[1'h0:1'h0];
  assign T4923 = T2943[1'h1:1'h1];
  assign T4924 = T4945 ? T4935 : T4925;
  assign T4925 = T4934 ? twiddle4_3_261_imag : twiddle4_3_260_imag;
  assign twiddle4_3_260_imag = T4928 + T4926;
  assign T4926 = $signed(T4927) / $signed(22'h100000);
  assign T4927 = $signed(31'h2b8ef77c) * $signed(16'hffff);
  assign T4928 = $signed(T4929) / $signed(22'h100000);
  assign T4929 = $signed(31'h511c3142) * $signed(16'h0);
  assign twiddle4_3_261_imag = T4932 + T4930;
  assign T4930 = $signed(T4931) / $signed(22'h100000);
  assign T4931 = $signed(31'h2b2003ab) * $signed(16'hffff);
  assign T4932 = $signed(T4933) / $signed(22'h100000);
  assign T4933 = $signed(31'h50b611f1) * $signed(16'h0);
  assign T4934 = T2943[1'h0:1'h0];
  assign T4935 = T4944 ? twiddle4_3_263_imag : twiddle4_3_262_imag;
  assign twiddle4_3_262_imag = T4938 + T4936;
  assign T4936 = $signed(T4937) / $signed(22'h100000);
  assign T4937 = $signed(31'h2ab02071) * $signed(16'hffff);
  assign T4938 = $signed(T4939) / $signed(22'h100000);
  assign T4939 = $signed(31'h5050f927) * $signed(16'h0);
  assign twiddle4_3_263_imag = T4942 + T4940;
  assign T4940 = $signed(T4941) / $signed(22'h100000);
  assign T4941 = $signed(31'h2a3f5039) * $signed(16'hffff);
  assign T4942 = $signed(T4943) / $signed(22'h100000);
  assign T4943 = $signed(31'h4fece916) * $signed(16'h0);
  assign T4944 = T2943[1'h0:1'h0];
  assign T4945 = T2943[1'h1:1'h1];
  assign T4946 = T2943[2'h2:2'h2];
  assign T4947 = T4992 ? T4970 : T4948;
  assign T4948 = T4969 ? T4959 : T4949;
  assign T4949 = T4958 ? twiddle4_3_265_imag : twiddle4_3_264_imag;
  assign twiddle4_3_264_imag = T4952 + T4950;
  assign T4950 = $signed(T4951) / $signed(22'h100000);
  assign T4951 = $signed(31'h29cd9577) * $signed(16'hffff);
  assign T4952 = $signed(T4953) / $signed(22'h100000);
  assign T4953 = $signed(31'h4f89e3e9) * $signed(16'h0);
  assign twiddle4_3_265_imag = T4956 + T4954;
  assign T4954 = $signed(T4955) / $signed(22'h100000);
  assign T4955 = $signed(31'h295af2a2) * $signed(16'hffff);
  assign T4956 = $signed(T4957) / $signed(22'h100000);
  assign T4957 = $signed(31'h4f27ebc5) * $signed(16'h0);
  assign T4958 = T2943[1'h0:1'h0];
  assign T4959 = T4968 ? twiddle4_3_267_imag : twiddle4_3_266_imag;
  assign twiddle4_3_266_imag = T4962 + T4960;
  assign T4960 = $signed(T4961) / $signed(22'h100000);
  assign T4961 = $signed(31'h28e76a37) * $signed(16'hffff);
  assign T4962 = $signed(T4963) / $signed(22'h100000);
  assign T4963 = $signed(31'h4ec702cc) * $signed(16'h0);
  assign twiddle4_3_267_imag = T4966 + T4964;
  assign T4964 = $signed(T4965) / $signed(22'h100000);
  assign T4965 = $signed(31'h2872feb6) * $signed(16'hffff);
  assign T4966 = $signed(T4967) / $signed(22'h100000);
  assign T4967 = $signed(31'h4e672b16) * $signed(16'h0);
  assign T4968 = T2943[1'h0:1'h0];
  assign T4969 = T2943[1'h1:1'h1];
  assign T4970 = T4991 ? T4981 : T4971;
  assign T4971 = T4980 ? twiddle4_3_269_imag : twiddle4_3_268_imag;
  assign twiddle4_3_268_imag = T4974 + T4972;
  assign T4972 = $signed(T4973) / $signed(22'h100000);
  assign T4973 = $signed(31'h27fdb2a6) * $signed(16'hffff);
  assign T4974 = $signed(T4975) / $signed(22'h100000);
  assign T4975 = $signed(31'h4e0866b9) * $signed(16'h0);
  assign twiddle4_3_269_imag = T4978 + T4976;
  assign T4976 = $signed(T4977) / $signed(22'h100000);
  assign T4977 = $signed(31'h27878893) * $signed(16'hffff);
  assign T4978 = $signed(T4979) / $signed(22'h100000);
  assign T4979 = $signed(31'h4daab7c1) * $signed(16'h0);
  assign T4980 = T2943[1'h0:1'h0];
  assign T4981 = T4990 ? twiddle4_3_271_imag : twiddle4_3_270_imag;
  assign twiddle4_3_270_imag = T4984 + T4982;
  assign T4982 = $signed(T4983) / $signed(22'h100000);
  assign T4983 = $signed(31'h2710830b) * $signed(16'hffff);
  assign T4984 = $signed(T4985) / $signed(22'h100000);
  assign T4985 = $signed(31'h4d4e2037) * $signed(16'h0);
  assign twiddle4_3_271_imag = T4988 + T4986;
  assign T4986 = $signed(T4987) / $signed(22'h100000);
  assign T4987 = $signed(31'h2698a4a5) * $signed(16'hffff);
  assign T4988 = $signed(T4989) / $signed(22'h100000);
  assign T4989 = $signed(31'h4cf2a21e) * $signed(16'h0);
  assign T4990 = T2943[1'h0:1'h0];
  assign T4991 = T2943[1'h1:1'h1];
  assign T4992 = T2943[2'h2:2'h2];
  assign T4993 = T2943[2'h3:2'h3];
  assign T4994 = T5093 ? T5041 : T4995;
  assign T4995 = T5040 ? T5018 : T4996;
  assign T4996 = T5017 ? T5007 : T4997;
  assign T4997 = T5006 ? twiddle4_3_273_imag : twiddle4_3_272_imag;
  assign twiddle4_3_272_imag = T5000 + T4998;
  assign T4998 = $signed(T4999) / $signed(22'h100000);
  assign T4999 = $signed(31'h261feff9) * $signed(16'hffff);
  assign T5000 = $signed(T5001) / $signed(22'h100000);
  assign T5001 = $signed(31'h4c983f71) * $signed(16'h0);
  assign twiddle4_3_273_imag = T5004 + T5002;
  assign T5002 = $signed(T5003) / $signed(22'h100000);
  assign T5003 = $signed(31'h25a667a6) * $signed(16'hffff);
  assign T5004 = $signed(T5005) / $signed(22'h100000);
  assign T5005 = $signed(31'h4c3efa25) * $signed(16'h0);
  assign T5006 = T2943[1'h0:1'h0];
  assign T5007 = T5016 ? twiddle4_3_275_imag : twiddle4_3_274_imag;
  assign twiddle4_3_274_imag = T5010 + T5008;
  assign T5008 = $signed(T5009) / $signed(22'h100000);
  assign T5009 = $signed(31'h252c0e4e) * $signed(16'hffff);
  assign T5010 = $signed(T5011) / $signed(22'h100000);
  assign T5011 = $signed(31'h4be6d42b) * $signed(16'h0);
  assign twiddle4_3_275_imag = T5014 + T5012;
  assign T5012 = $signed(T5013) / $signed(22'h100000);
  assign T5013 = $signed(31'h24b0e699) * $signed(16'hffff);
  assign T5014 = $signed(T5015) / $signed(22'h100000);
  assign T5015 = $signed(31'h4b8fcf6c) * $signed(16'h0);
  assign T5016 = T2943[1'h0:1'h0];
  assign T5017 = T2943[1'h1:1'h1];
  assign T5018 = T5039 ? T5029 : T5019;
  assign T5019 = T5028 ? twiddle4_3_277_imag : twiddle4_3_276_imag;
  assign twiddle4_3_276_imag = T5022 + T5020;
  assign T5020 = $signed(T5021) / $signed(22'h100000);
  assign T5021 = $signed(31'h2434f332) * $signed(16'hffff);
  assign T5022 = $signed(T5023) / $signed(22'h100000);
  assign T5023 = $signed(31'h4b39edca) * $signed(16'h0);
  assign twiddle4_3_277_imag = T5026 + T5024;
  assign T5024 = $signed(T5025) / $signed(22'h100000);
  assign T5025 = $signed(31'h23b836c9) * $signed(16'hffff);
  assign T5026 = $signed(T5027) / $signed(22'h100000);
  assign T5027 = $signed(31'h4ae53124) * $signed(16'h0);
  assign T5028 = T2943[1'h0:1'h0];
  assign T5029 = T5038 ? twiddle4_3_279_imag : twiddle4_3_278_imag;
  assign twiddle4_3_278_imag = T5032 + T5030;
  assign T5030 = $signed(T5031) / $signed(22'h100000);
  assign T5031 = $signed(31'h233ab413) * $signed(16'hffff);
  assign T5032 = $signed(T5033) / $signed(22'h100000);
  assign T5033 = $signed(31'h4a919b4e) * $signed(16'h0);
  assign twiddle4_3_279_imag = T5036 + T5034;
  assign T5034 = $signed(T5035) / $signed(22'h100000);
  assign T5035 = $signed(31'h22bc6dc9) * $signed(16'hffff);
  assign T5036 = $signed(T5037) / $signed(22'h100000);
  assign T5037 = $signed(31'h4a3f2e1a) * $signed(16'h0);
  assign T5038 = T2943[1'h0:1'h0];
  assign T5039 = T2943[1'h1:1'h1];
  assign T5040 = T2943[2'h2:2'h2];
  assign T5041 = T5092 ? T5064 : T5042;
  assign T5042 = T5063 ? T5053 : T5043;
  assign T5043 = T5052 ? twiddle4_3_281_imag : twiddle4_3_280_imag;
  assign twiddle4_3_280_imag = T5046 + T5044;
  assign T5044 = $signed(T5045) / $signed(22'h100000);
  assign T5045 = $signed(31'h223d66a8) * $signed(16'hffff);
  assign T5046 = $signed(T5047) / $signed(22'h100000);
  assign T5047 = $signed(31'h49edeb50) * $signed(16'h0);
  assign twiddle4_3_281_imag = T5050 + T5048;
  assign T5048 = $signed(T5049) / $signed(22'h100000);
  assign T5049 = $signed(31'h21bda170) * $signed(16'hffff);
  assign T5050 = $signed(T5051) / $signed(22'h100000);
  assign T5051 = $signed(31'h499dd4b5) * $signed(16'h0);
  assign T5052 = T2943[1'h0:1'h0];
  assign T5053 = T5062 ? twiddle4_3_283_imag : twiddle4_3_282_imag;
  assign twiddle4_3_282_imag = T5056 + T5054;
  assign T5054 = $signed(T5055) / $signed(22'h100000);
  assign T5055 = $signed(31'h213d20e8) * $signed(16'hffff);
  assign T5056 = $signed(T5057) / $signed(22'h100000);
  assign T5057 = $signed(31'h494eec03) * $signed(16'h0);
  assign twiddle4_3_283_imag = T5060 + T5058;
  assign T5058 = $signed(T5059) / $signed(22'h100000);
  assign T5059 = $signed(31'h20bbe7d8) * $signed(16'hffff);
  assign T5060 = $signed(T5061) / $signed(22'h100000);
  assign T5061 = $signed(31'h490132f3) * $signed(16'h0);
  assign T5062 = T2943[1'h0:1'h0];
  assign T5063 = T2943[1'h1:1'h1];
  assign T5064 = T5091 ? T5077 : T5065;
  assign T5065 = T5076 ? twiddle4_3_285_imag : twiddle4_3_284_imag;
  assign twiddle4_3_284_imag = T5068 + T5066;
  assign T5066 = $signed(T5067) / $signed(22'h100000);
  assign T5067 = $signed(31'h2039f90e) * $signed(16'hffff);
  assign T5068 = $signed(T5069) / $signed(22'h100000);
  assign T5069 = $signed(31'h48b4ab32) * $signed(16'h0);
  assign twiddle4_3_285_imag = T5074 + T5070;
  assign T5070 = {T5073, T5071};
  assign T5071 = $signed(T5072) / $signed(22'h100000);
  assign T5072 = $signed(30'h1fb7575c) * $signed(16'hffff);
  assign T5073 = T5071[6'h2d:6'h2d];
  assign T5074 = $signed(T5075) / $signed(22'h100000);
  assign T5075 = $signed(31'h4869566a) * $signed(16'h0);
  assign T5076 = T2943[1'h0:1'h0];
  assign T5077 = T5090 ? twiddle4_3_287_imag : twiddle4_3_286_imag;
  assign twiddle4_3_286_imag = T5082 + T5078;
  assign T5078 = {T5081, T5079};
  assign T5079 = $signed(T5080) / $signed(22'h100000);
  assign T5080 = $signed(30'h1f340596) * $signed(16'hffff);
  assign T5081 = T5079[6'h2d:6'h2d];
  assign T5082 = $signed(T5083) / $signed(22'h100000);
  assign T5083 = $signed(31'h481f363e) * $signed(16'h0);
  assign twiddle4_3_287_imag = T5088 + T5084;
  assign T5084 = {T5087, T5085};
  assign T5085 = $signed(T5086) / $signed(22'h100000);
  assign T5086 = $signed(30'h1eb00695) * $signed(16'hffff);
  assign T5087 = T5085[6'h2d:6'h2d];
  assign T5088 = $signed(T5089) / $signed(22'h100000);
  assign T5089 = $signed(31'h47d64c48) * $signed(16'h0);
  assign T5090 = T2943[1'h0:1'h0];
  assign T5091 = T2943[1'h1:1'h1];
  assign T5092 = T2943[2'h2:2'h2];
  assign T5093 = T2943[2'h3:2'h3];
  assign T5094 = T2943[3'h4:3'h4];
  assign T5095 = T5354 ? T5222 : T5096;
  assign T5096 = T5221 ? T5159 : T5097;
  assign T5097 = T5158 ? T5128 : T5098;
  assign T5098 = T5127 ? T5113 : T5099;
  assign T5099 = T5112 ? twiddle4_3_289_imag : twiddle4_3_288_imag;
  assign twiddle4_3_288_imag = T5104 + T5100;
  assign T5100 = {T5103, T5101};
  assign T5101 = $signed(T5102) / $signed(22'h100000);
  assign T5102 = $signed(30'h1e2b5d38) * $signed(16'hffff);
  assign T5103 = T5101[6'h2d:6'h2d];
  assign T5104 = $signed(T5105) / $signed(22'h100000);
  assign T5105 = $signed(31'h478e9a1d) * $signed(16'h0);
  assign twiddle4_3_289_imag = T5110 + T5106;
  assign T5106 = {T5109, T5107};
  assign T5107 = $signed(T5108) / $signed(22'h100000);
  assign T5108 = $signed(30'h1da60c5c) * $signed(16'hffff);
  assign T5109 = T5107[6'h2d:6'h2d];
  assign T5110 = $signed(T5111) / $signed(22'h100000);
  assign T5111 = $signed(31'h4748214d) * $signed(16'h0);
  assign T5112 = T2943[1'h0:1'h0];
  assign T5113 = T5126 ? twiddle4_3_291_imag : twiddle4_3_290_imag;
  assign twiddle4_3_290_imag = T5118 + T5114;
  assign T5114 = {T5117, T5115};
  assign T5115 = $signed(T5116) / $signed(22'h100000);
  assign T5116 = $signed(30'h1d2016e8) * $signed(16'hffff);
  assign T5117 = T5115[6'h2d:6'h2d];
  assign T5118 = $signed(T5119) / $signed(22'h100000);
  assign T5119 = $signed(31'h4702e35c) * $signed(16'h0);
  assign twiddle4_3_291_imag = T5124 + T5120;
  assign T5120 = {T5123, T5121};
  assign T5121 = $signed(T5122) / $signed(22'h100000);
  assign T5122 = $signed(30'h1c997fc3) * $signed(16'hffff);
  assign T5123 = T5121[6'h2d:6'h2d];
  assign T5124 = $signed(T5125) / $signed(22'h100000);
  assign T5125 = $signed(31'h46bee1cd) * $signed(16'h0);
  assign T5126 = T2943[1'h0:1'h0];
  assign T5127 = T2943[1'h1:1'h1];
  assign T5128 = T5157 ? T5143 : T5129;
  assign T5129 = T5142 ? twiddle4_3_293_imag : twiddle4_3_292_imag;
  assign twiddle4_3_292_imag = T5134 + T5130;
  assign T5130 = {T5133, T5131};
  assign T5131 = $signed(T5132) / $signed(22'h100000);
  assign T5132 = $signed(30'h1c1249d8) * $signed(16'hffff);
  assign T5133 = T5131[6'h2d:6'h2d];
  assign T5134 = $signed(T5135) / $signed(22'h100000);
  assign T5135 = $signed(31'h467c1e19) * $signed(16'h0);
  assign twiddle4_3_293_imag = T5140 + T5136;
  assign T5136 = {T5139, T5137};
  assign T5137 = $signed(T5138) / $signed(22'h100000);
  assign T5138 = $signed(30'h1b8a7814) * $signed(16'hffff);
  assign T5139 = T5137[6'h2d:6'h2d];
  assign T5140 = $signed(T5141) / $signed(22'h100000);
  assign T5141 = $signed(31'h463a99b1) * $signed(16'h0);
  assign T5142 = T2943[1'h0:1'h0];
  assign T5143 = T5156 ? twiddle4_3_295_imag : twiddle4_3_294_imag;
  assign twiddle4_3_294_imag = T5148 + T5144;
  assign T5144 = {T5147, T5145};
  assign T5145 = $signed(T5146) / $signed(22'h100000);
  assign T5146 = $signed(30'h1b020d6c) * $signed(16'hffff);
  assign T5147 = T5145[6'h2d:6'h2d];
  assign T5148 = $signed(T5149) / $signed(22'h100000);
  assign T5149 = $signed(31'h45fa5603) * $signed(16'h0);
  assign twiddle4_3_295_imag = T5154 + T5150;
  assign T5150 = {T5153, T5151};
  assign T5151 = $signed(T5152) / $signed(22'h100000);
  assign T5152 = $signed(30'h1a790cd3) * $signed(16'hffff);
  assign T5153 = T5151[6'h2d:6'h2d];
  assign T5154 = $signed(T5155) / $signed(22'h100000);
  assign T5155 = $signed(31'h45bb5473) * $signed(16'h0);
  assign T5156 = T2943[1'h0:1'h0];
  assign T5157 = T2943[1'h1:1'h1];
  assign T5158 = T2943[2'h2:2'h2];
  assign T5159 = T5220 ? T5190 : T5160;
  assign T5160 = T5189 ? T5175 : T5161;
  assign T5161 = T5174 ? twiddle4_3_297_imag : twiddle4_3_296_imag;
  assign twiddle4_3_296_imag = T5166 + T5162;
  assign T5162 = {T5165, T5163};
  assign T5163 = $signed(T5164) / $signed(22'h100000);
  assign T5164 = $signed(30'h19ef7943) * $signed(16'hffff);
  assign T5165 = T5163[6'h2d:6'h2d];
  assign T5166 = $signed(T5167) / $signed(22'h100000);
  assign T5167 = $signed(31'h457d965e) * $signed(16'h0);
  assign twiddle4_3_297_imag = T5172 + T5168;
  assign T5168 = {T5171, T5169};
  assign T5169 = $signed(T5170) / $signed(22'h100000);
  assign T5170 = $signed(30'h196555b7) * $signed(16'hffff);
  assign T5171 = T5169[6'h2d:6'h2d];
  assign T5172 = $signed(T5173) / $signed(22'h100000);
  assign T5173 = $signed(31'h45411d1b) * $signed(16'h0);
  assign T5174 = T2943[1'h0:1'h0];
  assign T5175 = T5188 ? twiddle4_3_299_imag : twiddle4_3_298_imag;
  assign twiddle4_3_298_imag = T5180 + T5176;
  assign T5176 = {T5179, T5177};
  assign T5177 = $signed(T5178) / $signed(22'h100000);
  assign T5178 = $signed(30'h18daa52e) * $signed(16'hffff);
  assign T5179 = T5177[6'h2d:6'h2d];
  assign T5180 = $signed(T5181) / $signed(22'h100000);
  assign T5181 = $signed(31'h4505e9fb) * $signed(16'h0);
  assign twiddle4_3_299_imag = T5186 + T5182;
  assign T5182 = {T5185, T5183};
  assign T5183 = $signed(T5184) / $signed(22'h100000);
  assign T5184 = $signed(30'h184f6aaa) * $signed(16'hffff);
  assign T5185 = T5183[6'h2d:6'h2d];
  assign T5186 = $signed(T5187) / $signed(22'h100000);
  assign T5187 = $signed(31'h44cbfe45) * $signed(16'h0);
  assign T5188 = T2943[1'h0:1'h0];
  assign T5189 = T2943[1'h1:1'h1];
  assign T5190 = T5219 ? T5205 : T5191;
  assign T5191 = T5204 ? twiddle4_3_301_imag : twiddle4_3_300_imag;
  assign twiddle4_3_300_imag = T5196 + T5192;
  assign T5192 = {T5195, T5193};
  assign T5193 = $signed(T5194) / $signed(22'h100000);
  assign T5194 = $signed(30'h17c3a931) * $signed(16'hffff);
  assign T5195 = T5193[6'h2d:6'h2d];
  assign T5196 = $signed(T5197) / $signed(22'h100000);
  assign T5197 = $signed(31'h44935b3c) * $signed(16'h0);
  assign twiddle4_3_301_imag = T5202 + T5198;
  assign T5198 = {T5201, T5199};
  assign T5199 = $signed(T5200) / $signed(22'h100000);
  assign T5200 = $signed(30'h173763c9) * $signed(16'hffff);
  assign T5201 = T5199[6'h2d:6'h2d];
  assign T5202 = $signed(T5203) / $signed(22'h100000);
  assign T5203 = $signed(31'h445c0219) * $signed(16'h0);
  assign T5204 = T2943[1'h0:1'h0];
  assign T5205 = T5218 ? twiddle4_3_303_imag : twiddle4_3_302_imag;
  assign twiddle4_3_302_imag = T5210 + T5206;
  assign T5206 = {T5209, T5207};
  assign T5207 = $signed(T5208) / $signed(22'h100000);
  assign T5208 = $signed(30'h16aa9d7d) * $signed(16'hffff);
  assign T5209 = T5207[6'h2d:6'h2d];
  assign T5210 = $signed(T5211) / $signed(22'h100000);
  assign T5211 = $signed(31'h4425f411) * $signed(16'h0);
  assign twiddle4_3_303_imag = T5216 + T5212;
  assign T5212 = {T5215, T5213};
  assign T5213 = $signed(T5214) / $signed(22'h100000);
  assign T5214 = $signed(30'h161d595c) * $signed(16'hffff);
  assign T5215 = T5213[6'h2d:6'h2d];
  assign T5216 = $signed(T5217) / $signed(22'h100000);
  assign T5217 = $signed(31'h43f1324e) * $signed(16'h0);
  assign T5218 = T2943[1'h0:1'h0];
  assign T5219 = T2943[1'h1:1'h1];
  assign T5220 = T2943[2'h2:2'h2];
  assign T5221 = T2943[2'h3:2'h3];
  assign T5222 = T5353 ? T5285 : T5223;
  assign T5223 = T5284 ? T5254 : T5224;
  assign T5224 = T5253 ? T5239 : T5225;
  assign T5225 = T5238 ? twiddle4_3_305_imag : twiddle4_3_304_imag;
  assign twiddle4_3_304_imag = T5230 + T5226;
  assign T5226 = {T5229, T5227};
  assign T5227 = $signed(T5228) / $signed(22'h100000);
  assign T5228 = $signed(30'h158f9a75) * $signed(16'hffff);
  assign T5229 = T5227[6'h2d:6'h2d];
  assign T5230 = $signed(T5231) / $signed(22'h100000);
  assign T5231 = $signed(31'h43bdbdf7) * $signed(16'h0);
  assign twiddle4_3_305_imag = T5236 + T5232;
  assign T5232 = {T5235, T5233};
  assign T5233 = $signed(T5234) / $signed(22'h100000);
  assign T5234 = $signed(30'h150163dc) * $signed(16'hffff);
  assign T5235 = T5233[6'h2d:6'h2d];
  assign T5236 = $signed(T5237) / $signed(22'h100000);
  assign T5237 = $signed(31'h438b9828) * $signed(16'h0);
  assign T5238 = T2943[1'h0:1'h0];
  assign T5239 = T5252 ? twiddle4_3_307_imag : twiddle4_3_306_imag;
  assign twiddle4_3_306_imag = T5244 + T5240;
  assign T5240 = {T5243, T5241};
  assign T5241 = $signed(T5242) / $signed(22'h100000);
  assign T5242 = $signed(30'h1472b8a5) * $signed(16'hffff);
  assign T5243 = T5241[6'h2d:6'h2d];
  assign T5244 = $signed(T5245) / $signed(22'h100000);
  assign T5245 = $signed(31'h435ac1f8) * $signed(16'h0);
  assign twiddle4_3_307_imag = T5250 + T5246;
  assign T5246 = {T5249, T5247};
  assign T5247 = $signed(T5248) / $signed(22'h100000);
  assign T5248 = $signed(30'h13e39be9) * $signed(16'hffff);
  assign T5249 = T5247[6'h2d:6'h2d];
  assign T5250 = $signed(T5251) / $signed(22'h100000);
  assign T5251 = $signed(31'h432b3c76) * $signed(16'h0);
  assign T5252 = T2943[1'h0:1'h0];
  assign T5253 = T2943[1'h1:1'h1];
  assign T5254 = T5283 ? T5269 : T5255;
  assign T5255 = T5268 ? twiddle4_3_309_imag : twiddle4_3_308_imag;
  assign twiddle4_3_308_imag = T5260 + T5256;
  assign T5256 = {T5259, T5257};
  assign T5257 = $signed(T5258) / $signed(22'h100000);
  assign T5258 = $signed(30'h135410c2) * $signed(16'hffff);
  assign T5259 = T5257[6'h2d:6'h2d];
  assign T5260 = $signed(T5261) / $signed(22'h100000);
  assign T5261 = $signed(31'h42fd08aa) * $signed(16'h0);
  assign twiddle4_3_309_imag = T5266 + T5262;
  assign T5262 = {T5265, T5263};
  assign T5263 = $signed(T5264) / $signed(22'h100000);
  assign T5264 = $signed(30'h12c41a4e) * $signed(16'hffff);
  assign T5265 = T5263[6'h2d:6'h2d];
  assign T5266 = $signed(T5267) / $signed(22'h100000);
  assign T5267 = $signed(31'h42d02794) * $signed(16'h0);
  assign T5268 = T2943[1'h0:1'h0];
  assign T5269 = T5282 ? twiddle4_3_311_imag : twiddle4_3_310_imag;
  assign twiddle4_3_310_imag = T5274 + T5270;
  assign T5270 = {T5273, T5271};
  assign T5271 = $signed(T5272) / $signed(22'h100000);
  assign T5272 = $signed(30'h1233bbab) * $signed(16'hffff);
  assign T5273 = T5271[6'h2d:6'h2d];
  assign T5274 = $signed(T5275) / $signed(22'h100000);
  assign T5275 = $signed(31'h42a49a2f) * $signed(16'h0);
  assign twiddle4_3_311_imag = T5280 + T5276;
  assign T5276 = {T5279, T5277};
  assign T5277 = $signed(T5278) / $signed(22'h100000);
  assign T5278 = $signed(30'h11a2f7fb) * $signed(16'hffff);
  assign T5279 = T5277[6'h2d:6'h2d];
  assign T5280 = $signed(T5281) / $signed(22'h100000);
  assign T5281 = $signed(31'h427a616a) * $signed(16'h0);
  assign T5282 = T2943[1'h0:1'h0];
  assign T5283 = T2943[1'h1:1'h1];
  assign T5284 = T2943[2'h2:2'h2];
  assign T5285 = T5352 ? T5318 : T5286;
  assign T5286 = T5317 ? T5301 : T5287;
  assign T5287 = T5300 ? twiddle4_3_313_imag : twiddle4_3_312_imag;
  assign twiddle4_3_312_imag = T5292 + T5288;
  assign T5288 = {T5291, T5289};
  assign T5289 = $signed(T5290) / $signed(22'h100000);
  assign T5290 = $signed(30'h1111d262) * $signed(16'hffff);
  assign T5291 = T5289[6'h2d:6'h2d];
  assign T5292 = $signed(T5293) / $signed(22'h100000);
  assign T5293 = $signed(31'h42517e32) * $signed(16'h0);
  assign twiddle4_3_313_imag = T5298 + T5294;
  assign T5294 = {T5297, T5295};
  assign T5295 = $signed(T5296) / $signed(22'h100000);
  assign T5296 = $signed(30'h10804e05) * $signed(16'hffff);
  assign T5297 = T5295[6'h2d:6'h2d];
  assign T5298 = $signed(T5299) / $signed(22'h100000);
  assign T5299 = $signed(31'h4229f168) * $signed(16'h0);
  assign T5300 = T2943[1'h0:1'h0];
  assign T5301 = T5316 ? twiddle4_3_315_imag : twiddle4_3_314_imag;
  assign twiddle4_3_314_imag = T5307 + T5302;
  assign T5302 = {T5305, T5303};
  assign T5303 = $signed(T5304) / $signed(22'h100000);
  assign T5304 = $signed(29'hfee6e0d) * $signed(16'hffff);
  assign T5305 = T5306 ? 2'h3 : 2'h0;
  assign T5306 = T5303[6'h2c:6'h2c];
  assign T5307 = $signed(T5308) / $signed(22'h100000);
  assign T5308 = $signed(31'h4203bbe8) * $signed(16'h0);
  assign twiddle4_3_315_imag = T5314 + T5309;
  assign T5309 = {T5312, T5310};
  assign T5310 = $signed(T5311) / $signed(22'h100000);
  assign T5311 = $signed(29'hf5c35a3) * $signed(16'hffff);
  assign T5312 = T5313 ? 2'h3 : 2'h0;
  assign T5313 = T5310[6'h2c:6'h2c];
  assign T5314 = $signed(T5315) / $signed(22'h100000);
  assign T5315 = $signed(31'h41dede87) * $signed(16'h0);
  assign T5316 = T2943[1'h0:1'h0];
  assign T5317 = T2943[1'h1:1'h1];
  assign T5318 = T5351 ? T5335 : T5319;
  assign T5319 = T5334 ? twiddle4_3_317_imag : twiddle4_3_316_imag;
  assign twiddle4_3_316_imag = T5325 + T5320;
  assign T5320 = {T5323, T5321};
  assign T5321 = $signed(T5322) / $signed(22'h100000);
  assign T5322 = $signed(29'hec9a7f2) * $signed(16'hffff);
  assign T5323 = T5324 ? 2'h3 : 2'h0;
  assign T5324 = T5321[6'h2c:6'h2c];
  assign T5325 = $signed(T5326) / $signed(22'h100000);
  assign T5326 = $signed(31'h41bb5a12) * $signed(16'h0);
  assign twiddle4_3_317_imag = T5332 + T5327;
  assign T5327 = {T5330, T5328};
  assign T5328 = $signed(T5329) / $signed(22'h100000);
  assign T5329 = $signed(29'he36c829) * $signed(16'hffff);
  assign T5330 = T5331 ? 2'h3 : 2'h0;
  assign T5331 = T5328[6'h2c:6'h2c];
  assign T5332 = $signed(T5333) / $signed(22'h100000);
  assign T5333 = $signed(31'h41992f4c) * $signed(16'h0);
  assign T5334 = T2943[1'h0:1'h0];
  assign T5335 = T5350 ? twiddle4_3_319_imag : twiddle4_3_318_imag;
  assign twiddle4_3_318_imag = T5341 + T5336;
  assign T5336 = {T5339, T5337};
  assign T5337 = $signed(T5338) / $signed(22'h100000);
  assign T5338 = $signed(29'hda39977) * $signed(16'hffff);
  assign T5339 = T5340 ? 2'h3 : 2'h0;
  assign T5340 = T5337[6'h2c:6'h2c];
  assign T5341 = $signed(T5342) / $signed(22'h100000);
  assign T5342 = $signed(31'h41785ef5) * $signed(16'h0);
  assign twiddle4_3_319_imag = T5348 + T5343;
  assign T5343 = {T5346, T5344};
  assign T5344 = $signed(T5345) / $signed(22'h100000);
  assign T5345 = $signed(29'hd101f0d) * $signed(16'hffff);
  assign T5346 = T5347 ? 2'h3 : 2'h0;
  assign T5347 = T5344[6'h2c:6'h2c];
  assign T5348 = $signed(T5349) / $signed(22'h100000);
  assign T5349 = $signed(31'h4158e9c1) * $signed(16'h0);
  assign T5350 = T2943[1'h0:1'h0];
  assign T5351 = T2943[1'h1:1'h1];
  assign T5352 = T2943[2'h2:2'h2];
  assign T5353 = T2943[2'h3:2'h3];
  assign T5354 = T2943[3'h4:3'h4];
  assign T5355 = T2943[3'h5:3'h5];
  assign T5356 = T5914 ? T5643 : T5357;
  assign T5357 = T5642 ? T5500 : T5358;
  assign T5358 = T5499 ? T5429 : T5359;
  assign T5359 = T5428 ? T5394 : T5360;
  assign T5360 = T5393 ? T5377 : T5361;
  assign T5361 = T5376 ? twiddle4_3_321_imag : twiddle4_3_320_imag;
  assign twiddle4_3_320_imag = T5367 + T5362;
  assign T5362 = {T5365, T5363};
  assign T5363 = $signed(T5364) / $signed(22'h100000);
  assign T5364 = $signed(29'hc7c5c1e) * $signed(16'hffff);
  assign T5365 = T5366 ? 2'h3 : 2'h0;
  assign T5366 = T5363[6'h2c:6'h2c];
  assign T5367 = $signed(T5368) / $signed(22'h100000);
  assign T5368 = $signed(31'h413ad061) * $signed(16'h0);
  assign twiddle4_3_321_imag = T5374 + T5369;
  assign T5369 = {T5372, T5370};
  assign T5370 = $signed(T5371) / $signed(22'h100000);
  assign T5371 = $signed(29'hbe853dd) * $signed(16'hffff);
  assign T5372 = T5373 ? 2'h3 : 2'h0;
  assign T5373 = T5370[6'h2c:6'h2c];
  assign T5374 = $signed(T5375) / $signed(22'h100000);
  assign T5375 = $signed(31'h411e137a) * $signed(16'h0);
  assign T5376 = T2943[1'h0:1'h0];
  assign T5377 = T5392 ? twiddle4_3_323_imag : twiddle4_3_322_imag;
  assign twiddle4_3_322_imag = T5383 + T5378;
  assign T5378 = {T5381, T5379};
  assign T5379 = $signed(T5380) / $signed(22'h100000);
  assign T5380 = $signed(29'hb540982) * $signed(16'hffff);
  assign T5381 = T5382 ? 2'h3 : 2'h0;
  assign T5382 = T5379[6'h2c:6'h2c];
  assign T5383 = $signed(T5384) / $signed(22'h100000);
  assign T5384 = $signed(31'h4102b3ad) * $signed(16'h0);
  assign twiddle4_3_323_imag = T5390 + T5385;
  assign T5385 = {T5388, T5386};
  assign T5386 = $signed(T5387) / $signed(22'h100000);
  assign T5387 = $signed(29'habf8043) * $signed(16'hffff);
  assign T5388 = T5389 ? 2'h3 : 2'h0;
  assign T5389 = T5386[6'h2c:6'h2c];
  assign T5390 = $signed(T5391) / $signed(22'h100000);
  assign T5391 = $signed(31'h40e8b191) * $signed(16'h0);
  assign T5392 = T2943[1'h0:1'h0];
  assign T5393 = T2943[1'h1:1'h1];
  assign T5394 = T5427 ? T5411 : T5395;
  assign T5395 = T5410 ? twiddle4_3_325_imag : twiddle4_3_324_imag;
  assign twiddle4_3_324_imag = T5401 + T5396;
  assign T5396 = {T5399, T5397};
  assign T5397 = $signed(T5398) / $signed(22'h100000);
  assign T5398 = $signed(29'ha2abb58) * $signed(16'hffff);
  assign T5399 = T5400 ? 2'h3 : 2'h0;
  assign T5400 = T5397[6'h2c:6'h2c];
  assign T5401 = $signed(T5402) / $signed(22'h100000);
  assign T5402 = $signed(31'h40d00db7) * $signed(16'h0);
  assign twiddle4_3_325_imag = T5408 + T5403;
  assign T5403 = {T5406, T5404};
  assign T5404 = $signed(T5405) / $signed(22'h100000);
  assign T5405 = $signed(29'h995bdfc) * $signed(16'hffff);
  assign T5406 = T5407 ? 2'h3 : 2'h0;
  assign T5407 = T5404[6'h2c:6'h2c];
  assign T5408 = $signed(T5409) / $signed(22'h100000);
  assign T5409 = $signed(31'h40b8c8a8) * $signed(16'h0);
  assign T5410 = T2943[1'h0:1'h0];
  assign T5411 = T5426 ? twiddle4_3_327_imag : twiddle4_3_326_imag;
  assign twiddle4_3_326_imag = T5417 + T5412;
  assign T5412 = {T5415, T5413};
  assign T5413 = $signed(T5414) / $signed(22'h100000);
  assign T5414 = $signed(29'h9008b6a) * $signed(16'hffff);
  assign T5415 = T5416 ? 2'h3 : 2'h0;
  assign T5416 = T5413[6'h2c:6'h2c];
  assign T5417 = $signed(T5418) / $signed(22'h100000);
  assign T5418 = $signed(31'h40a2e2e4) * $signed(16'h0);
  assign twiddle4_3_327_imag = T5424 + T5419;
  assign T5419 = {T5422, T5420};
  assign T5420 = $signed(T5421) / $signed(22'h100000);
  assign T5421 = $signed(29'h86b26de) * $signed(16'hffff);
  assign T5422 = T5423 ? 2'h3 : 2'h0;
  assign T5423 = T5420[6'h2c:6'h2c];
  assign T5424 = $signed(T5425) / $signed(22'h100000);
  assign T5425 = $signed(31'h408e5ce6) * $signed(16'h0);
  assign T5426 = T2943[1'h0:1'h0];
  assign T5427 = T2943[1'h1:1'h1];
  assign T5428 = T2943[2'h2:2'h2];
  assign T5429 = T5498 ? T5464 : T5430;
  assign T5430 = T5463 ? T5447 : T5431;
  assign T5431 = T5446 ? twiddle4_3_329_imag : twiddle4_3_328_imag;
  assign twiddle4_3_328_imag = T5437 + T5432;
  assign T5432 = {T5435, T5433};
  assign T5433 = $signed(T5434) / $signed(22'h100000);
  assign T5434 = $signed(28'h7d59395) * $signed(16'hffff);
  assign T5435 = T5436 ? 3'h7 : 3'h0;
  assign T5436 = T5433[6'h2b:6'h2b];
  assign T5437 = $signed(T5438) / $signed(22'h100000);
  assign T5438 = $signed(31'h407b371f) * $signed(16'h0);
  assign twiddle4_3_329_imag = T5444 + T5439;
  assign T5439 = {T5442, T5440};
  assign T5440 = $signed(T5441) / $signed(22'h100000);
  assign T5441 = $signed(28'h73fd4ce) * $signed(16'hffff);
  assign T5442 = T5443 ? 3'h7 : 3'h0;
  assign T5443 = T5440[6'h2b:6'h2b];
  assign T5444 = $signed(T5445) / $signed(22'h100000);
  assign T5445 = $signed(31'h406971f9) * $signed(16'h0);
  assign T5446 = T2943[1'h0:1'h0];
  assign T5447 = T5462 ? twiddle4_3_331_imag : twiddle4_3_330_imag;
  assign twiddle4_3_330_imag = T5453 + T5448;
  assign T5448 = {T5451, T5449};
  assign T5449 = $signed(T5450) / $signed(22'h100000);
  assign T5450 = $signed(28'h6a9edc9) * $signed(16'hffff);
  assign T5451 = T5452 ? 3'h7 : 3'h0;
  assign T5452 = T5449[6'h2b:6'h2b];
  assign T5453 = $signed(T5454) / $signed(22'h100000);
  assign T5454 = $signed(31'h40590dd8) * $signed(16'h0);
  assign twiddle4_3_331_imag = T5460 + T5455;
  assign T5455 = {T5458, T5456};
  assign T5456 = $signed(T5457) / $signed(22'h100000);
  assign T5457 = $signed(28'h613e1c4) * $signed(16'hffff);
  assign T5458 = T5459 ? 3'h7 : 3'h0;
  assign T5459 = T5456[6'h2b:6'h2b];
  assign T5460 = $signed(T5461) / $signed(22'h100000);
  assign T5461 = $signed(31'h404a0b16) * $signed(16'h0);
  assign T5462 = T2943[1'h0:1'h0];
  assign T5463 = T2943[1'h1:1'h1];
  assign T5464 = T5497 ? T5481 : T5465;
  assign T5465 = T5480 ? twiddle4_3_333_imag : twiddle4_3_332_imag;
  assign twiddle4_3_332_imag = T5471 + T5466;
  assign T5466 = {T5469, T5467};
  assign T5467 = $signed(T5468) / $signed(22'h100000);
  assign T5468 = $signed(28'h57db402) * $signed(16'hffff);
  assign T5469 = T5470 ? 3'h7 : 3'h0;
  assign T5470 = T5467[6'h2b:6'h2b];
  assign T5471 = $signed(T5472) / $signed(22'h100000);
  assign T5472 = $signed(31'h403c6a07) * $signed(16'h0);
  assign twiddle4_3_333_imag = T5478 + T5473;
  assign T5473 = {T5476, T5474};
  assign T5474 = $signed(T5475) / $signed(22'h100000);
  assign T5475 = $signed(28'h4e767c4) * $signed(16'hffff);
  assign T5476 = T5477 ? 3'h7 : 3'h0;
  assign T5477 = T5474[6'h2b:6'h2b];
  assign T5478 = $signed(T5479) / $signed(22'h100000);
  assign T5479 = $signed(31'h40302af6) * $signed(16'h0);
  assign T5480 = T2943[1'h0:1'h0];
  assign T5481 = T5496 ? twiddle4_3_335_imag : twiddle4_3_334_imag;
  assign twiddle4_3_334_imag = T5487 + T5482;
  assign T5482 = {T5485, T5483};
  assign T5483 = $signed(T5484) / $signed(22'h100000);
  assign T5484 = $signed(28'h451004d) * $signed(16'hffff);
  assign T5485 = T5486 ? 3'h7 : 3'h0;
  assign T5486 = T5483[6'h2b:6'h2b];
  assign T5487 = $signed(T5488) / $signed(22'h100000);
  assign T5488 = $signed(31'h40254e27) * $signed(16'h0);
  assign twiddle4_3_335_imag = T5494 + T5489;
  assign T5489 = {T5492, T5490};
  assign T5490 = $signed(T5491) / $signed(22'h100000);
  assign T5491 = $signed(27'h3ba80df) * $signed(16'hffff);
  assign T5492 = T5493 ? 4'hf : 4'h0;
  assign T5493 = T5490[6'h2a:6'h2a];
  assign T5494 = $signed(T5495) / $signed(22'h100000);
  assign T5495 = $signed(31'h401bd3d7) * $signed(16'h0);
  assign T5496 = T2943[1'h0:1'h0];
  assign T5497 = T2943[1'h1:1'h1];
  assign T5498 = T2943[2'h2:2'h2];
  assign T5499 = T2943[2'h3:2'h3];
  assign T5500 = T5641 ? T5571 : T5501;
  assign T5501 = T5570 ? T5536 : T5502;
  assign T5502 = T5535 ? T5519 : T5503;
  assign T5503 = T5518 ? twiddle4_3_337_imag : twiddle4_3_336_imag;
  assign twiddle4_3_336_imag = T5509 + T5504;
  assign T5504 = {T5507, T5505};
  assign T5505 = $signed(T5506) / $signed(22'h100000);
  assign T5506 = $signed(27'h323ecbe) * $signed(16'hffff);
  assign T5507 = T5508 ? 4'hf : 4'h0;
  assign T5508 = T5505[6'h2a:6'h2a];
  assign T5509 = $signed(T5510) / $signed(22'h100000);
  assign T5510 = $signed(31'h4013bc3a) * $signed(16'h0);
  assign twiddle4_3_337_imag = T5516 + T5511;
  assign T5511 = {T5514, T5512};
  assign T5512 = $signed(T5513) / $signed(22'h100000);
  assign T5513 = $signed(27'h28d472d) * $signed(16'hffff);
  assign T5514 = T5515 ? 4'hf : 4'h0;
  assign T5515 = T5512[6'h2a:6'h2a];
  assign T5516 = $signed(T5517) / $signed(22'h100000);
  assign T5517 = $signed(31'h400d077c) * $signed(16'h0);
  assign T5518 = T2943[1'h0:1'h0];
  assign T5519 = T5534 ? twiddle4_3_339_imag : twiddle4_3_338_imag;
  assign twiddle4_3_338_imag = T5525 + T5520;
  assign T5520 = {T5523, T5521};
  assign T5521 = $signed(T5522) / $signed(22'h100000);
  assign T5522 = $signed(26'h1f69373) * $signed(16'hffff);
  assign T5523 = T5524 ? 5'h1f : 5'h0;
  assign T5524 = T5521[6'h29:6'h29];
  assign T5525 = $signed(T5526) / $signed(22'h100000);
  assign T5526 = $signed(31'h4007b5c5) * $signed(16'h0);
  assign twiddle4_3_339_imag = T5532 + T5527;
  assign T5527 = {T5530, T5528};
  assign T5528 = $signed(T5529) / $signed(22'h100000);
  assign T5529 = $signed(26'h15fd4d2) * $signed(16'hffff);
  assign T5530 = T5531 ? 5'h1f : 5'h0;
  assign T5531 = T5528[6'h29:6'h29];
  assign T5532 = $signed(T5533) / $signed(22'h100000);
  assign T5533 = $signed(31'h4003c730) * $signed(16'h0);
  assign T5534 = T2943[1'h0:1'h0];
  assign T5535 = T2943[1'h1:1'h1];
  assign T5536 = T5569 ? T5553 : T5537;
  assign T5537 = T5552 ? twiddle4_3_341_imag : twiddle4_3_340_imag;
  assign twiddle4_3_340_imag = T5543 + T5538;
  assign T5538 = {T5541, T5539};
  assign T5539 = $signed(T5540) / $signed(22'h100000);
  assign T5540 = $signed(25'hc90e8f) * $signed(16'hffff);
  assign T5541 = T5542 ? 6'h3f : 6'h0;
  assign T5542 = T5539[6'h28:6'h28];
  assign T5543 = $signed(T5544) / $signed(22'h100000);
  assign T5544 = $signed(31'h40013bd3) * $signed(16'h0);
  assign twiddle4_3_341_imag = T5550 + T5545;
  assign T5545 = {T5548, T5546};
  assign T5546 = $signed(T5547) / $signed(22'h100000);
  assign T5547 = $signed(23'h3243f1) * $signed(16'hffff);
  assign T5548 = T5549 ? 8'hff : 8'h0;
  assign T5549 = T5546[6'h26:6'h26];
  assign T5550 = $signed(T5551) / $signed(22'h100000);
  assign T5551 = $signed(31'h400013be) * $signed(16'h0);
  assign T5552 = T2943[1'h0:1'h0];
  assign T5553 = T5568 ? twiddle4_3_343_imag : twiddle4_3_342_imag;
  assign twiddle4_3_342_imag = T5559 + T5554;
  assign T5554 = {T5557, T5555};
  assign T5555 = $signed(T5556) / $signed(22'h100000);
  assign T5556 = $signed(24'h9b783d) * $signed(16'hffff);
  assign T5557 = T5558 ? 7'h7f : 7'h0;
  assign T5558 = T5555[6'h27:6'h27];
  assign T5559 = $signed(T5560) / $signed(22'h100000);
  assign T5560 = $signed(31'h40004ef5) * $signed(16'h0);
  assign twiddle4_3_343_imag = T5566 + T5561;
  assign T5561 = {T5564, T5562};
  assign T5562 = $signed(T5563) / $signed(22'h100000);
  assign T5563 = $signed(25'h104aeb5) * $signed(16'hffff);
  assign T5564 = T5565 ? 6'h3f : 6'h0;
  assign T5565 = T5562[6'h28:6'h28];
  assign T5566 = $signed(T5567) / $signed(22'h100000);
  assign T5567 = $signed(31'h4001ed79) * $signed(16'h0);
  assign T5568 = T2943[1'h0:1'h0];
  assign T5569 = T2943[1'h1:1'h1];
  assign T5570 = T2943[2'h2:2'h2];
  assign T5571 = T5640 ? T5606 : T5572;
  assign T5572 = T5605 ? T5589 : T5573;
  assign T5573 = T5588 ? twiddle4_3_345_imag : twiddle4_3_344_imag;
  assign twiddle4_3_344_imag = T5579 + T5574;
  assign T5574 = {T5577, T5575};
  assign T5575 = $signed(T5576) / $signed(22'h100000);
  assign T5576 = $signed(26'h26deaa1) * $signed(16'hffff);
  assign T5577 = T5578 ? 5'h1f : 5'h0;
  assign T5578 = T5575[6'h29:6'h29];
  assign T5579 = $signed(T5580) / $signed(22'h100000);
  assign T5580 = $signed(31'h4004ef3f) * $signed(16'h0);
  assign twiddle4_3_345_imag = T5586 + T5581;
  assign T5581 = {T5584, T5582};
  assign T5582 = $signed(T5583) / $signed(22'h100000);
  assign T5583 = $signed(27'h5d72f45) * $signed(16'hffff);
  assign T5584 = T5585 ? 4'hf : 4'h0;
  assign T5585 = T5582[6'h2a:6'h2a];
  assign T5586 = $signed(T5587) / $signed(22'h100000);
  assign T5587 = $signed(31'h40095438) * $signed(16'h0);
  assign T5588 = T2943[1'h0:1'h0];
  assign T5589 = T5604 ? twiddle4_3_347_imag : twiddle4_3_346_imag;
  assign twiddle4_3_346_imag = T5595 + T5590;
  assign T5590 = {T5593, T5591};
  assign T5591 = $signed(T5592) / $signed(22'h100000);
  assign T5592 = $signed(27'h5407fe6) * $signed(16'hffff);
  assign T5593 = T5594 ? 4'hf : 4'h0;
  assign T5594 = T5591[6'h2a:6'h2a];
  assign T5595 = $signed(T5596) / $signed(22'h100000);
  assign T5596 = $signed(31'h400f1c4b) * $signed(16'h0);
  assign twiddle4_3_347_imag = T5602 + T5597;
  assign T5597 = {T5600, T5598};
  assign T5598 = $signed(T5599) / $signed(22'h100000);
  assign T5599 = $signed(27'h4a9dfc9) * $signed(16'hffff);
  assign T5600 = T5601 ? 4'hf : 4'h0;
  assign T5601 = T5598[6'h2a:6'h2a];
  assign T5602 = $signed(T5603) / $signed(22'h100000);
  assign T5603 = $signed(31'h40164757) * $signed(16'h0);
  assign T5604 = T2943[1'h0:1'h0];
  assign T5605 = T2943[1'h1:1'h1];
  assign T5606 = T5639 ? T5623 : T5607;
  assign T5607 = T5622 ? twiddle4_3_349_imag : twiddle4_3_348_imag;
  assign twiddle4_3_348_imag = T5613 + T5608;
  assign T5608 = {T5611, T5609};
  assign T5609 = $signed(T5610) / $signed(22'h100000);
  assign T5610 = $signed(27'h4135231) * $signed(16'hffff);
  assign T5611 = T5612 ? 4'hf : 4'h0;
  assign T5612 = T5609[6'h2a:6'h2a];
  assign T5613 = $signed(T5614) / $signed(22'h100000);
  assign T5614 = $signed(31'h401ed535) * $signed(16'h0);
  assign twiddle4_3_349_imag = T5620 + T5615;
  assign T5615 = {T5618, T5616};
  assign T5616 = $signed(T5617) / $signed(22'h100000);
  assign T5617 = $signed(28'hb7cda63) * $signed(16'hffff);
  assign T5618 = T5619 ? 3'h7 : 3'h0;
  assign T5619 = T5616[6'h2b:6'h2b];
  assign T5620 = $signed(T5621) / $signed(22'h100000);
  assign T5621 = $signed(31'h4028c5b6) * $signed(16'h0);
  assign T5622 = T2943[1'h0:1'h0];
  assign T5623 = T5638 ? twiddle4_3_351_imag : twiddle4_3_350_imag;
  assign twiddle4_3_350_imag = T5629 + T5624;
  assign T5624 = {T5627, T5625};
  assign T5625 = $signed(T5626) / $signed(22'h100000);
  assign T5626 = $signed(28'hae67ba2) * $signed(16'hffff);
  assign T5627 = T5628 ? 3'h7 : 3'h0;
  assign T5628 = T5625[6'h2b:6'h2b];
  assign T5629 = $signed(T5630) / $signed(22'h100000);
  assign T5630 = $signed(31'h403418a2) * $signed(16'h0);
  assign twiddle4_3_351_imag = T5636 + T5631;
  assign T5631 = {T5634, T5632};
  assign T5632 = $signed(T5633) / $signed(22'h100000);
  assign T5633 = $signed(28'ha503931) * $signed(16'hffff);
  assign T5634 = T5635 ? 3'h7 : 3'h0;
  assign T5635 = T5632[6'h2b:6'h2b];
  assign T5636 = $signed(T5637) / $signed(22'h100000);
  assign T5637 = $signed(31'h4040cdbb) * $signed(16'h0);
  assign T5638 = T2943[1'h0:1'h0];
  assign T5639 = T2943[1'h1:1'h1];
  assign T5640 = T2943[2'h2:2'h2];
  assign T5641 = T2943[2'h3:2'h3];
  assign T5642 = T2943[3'h4:3'h4];
  assign T5643 = T5913 ? T5786 : T5644;
  assign T5644 = T5785 ? T5715 : T5645;
  assign T5645 = T5714 ? T5680 : T5646;
  assign T5646 = T5679 ? T5663 : T5647;
  assign T5647 = T5662 ? twiddle4_3_353_imag : twiddle4_3_352_imag;
  assign twiddle4_3_352_imag = T5653 + T5648;
  assign T5648 = {T5651, T5649};
  assign T5649 = $signed(T5650) / $signed(22'h100000);
  assign T5650 = $signed(28'h9ba1651) * $signed(16'hffff);
  assign T5651 = T5652 ? 3'h7 : 3'h0;
  assign T5652 = T5649[6'h2b:6'h2b];
  assign T5653 = $signed(T5654) / $signed(22'h100000);
  assign T5654 = $signed(31'h404ee4b9) * $signed(16'h0);
  assign twiddle4_3_353_imag = T5660 + T5655;
  assign T5655 = {T5658, T5656};
  assign T5656 = $signed(T5657) / $signed(22'h100000);
  assign T5657 = $signed(28'h9241645) * $signed(16'hffff);
  assign T5658 = T5659 ? 3'h7 : 3'h0;
  assign T5659 = T5656[6'h2b:6'h2b];
  assign T5660 = $signed(T5661) / $signed(22'h100000);
  assign T5661 = $signed(31'h405e5d4f) * $signed(16'h0);
  assign T5662 = T2943[1'h0:1'h0];
  assign T5663 = T5678 ? twiddle4_3_355_imag : twiddle4_3_354_imag;
  assign twiddle4_3_354_imag = T5669 + T5664;
  assign T5664 = {T5667, T5665};
  assign T5665 = $signed(T5666) / $signed(22'h100000);
  assign T5666 = $signed(28'h88e3c4e) * $signed(16'hffff);
  assign T5667 = T5668 ? 3'h7 : 3'h0;
  assign T5668 = T5665[6'h2b:6'h2b];
  assign T5669 = $signed(T5670) / $signed(22'h100000);
  assign T5670 = $signed(31'h406f3727) * $signed(16'h0);
  assign twiddle4_3_355_imag = T5676 + T5671;
  assign T5671 = {T5674, T5672};
  assign T5672 = $signed(T5673) / $signed(22'h100000);
  assign T5673 = $signed(29'h17f88baa) * $signed(16'hffff);
  assign T5674 = T5675 ? 2'h3 : 2'h0;
  assign T5675 = T5672[6'h2c:6'h2c];
  assign T5676 = $signed(T5677) / $signed(22'h100000);
  assign T5677 = $signed(31'h408171e2) * $signed(16'h0);
  assign T5678 = T2943[1'h0:1'h0];
  assign T5679 = T2943[1'h1:1'h1];
  assign T5680 = T5713 ? T5697 : T5681;
  assign T5681 = T5696 ? twiddle4_3_357_imag : twiddle4_3_356_imag;
  assign twiddle4_3_356_imag = T5687 + T5682;
  assign T5682 = {T5685, T5683};
  assign T5683 = $signed(T5684) / $signed(22'h100000);
  assign T5684 = $signed(29'h17630799) * $signed(16'hffff);
  assign T5685 = T5686 ? 2'h3 : 2'h0;
  assign T5686 = T5683[6'h2c:6'h2c];
  assign T5687 = $signed(T5688) / $signed(22'h100000);
  assign T5688 = $signed(31'h40950d1d) * $signed(16'h0);
  assign twiddle4_3_357_imag = T5694 + T5689;
  assign T5689 = {T5692, T5690};
  assign T5690 = $signed(T5691) / $signed(22'h100000);
  assign T5691 = $signed(29'h16cdb35a) * $signed(16'hffff);
  assign T5692 = T5693 ? 2'h3 : 2'h0;
  assign T5693 = T5690[6'h2c:6'h2c];
  assign T5694 = $signed(T5695) / $signed(22'h100000);
  assign T5695 = $signed(31'h40aa086a) * $signed(16'h0);
  assign T5696 = T2943[1'h0:1'h0];
  assign T5697 = T5712 ? twiddle4_3_359_imag : twiddle4_3_358_imag;
  assign twiddle4_3_358_imag = T5703 + T5698;
  assign T5698 = {T5701, T5699};
  assign T5699 = $signed(T5700) / $signed(22'h100000);
  assign T5700 = $signed(29'h16389228) * $signed(16'hffff);
  assign T5701 = T5702 ? 2'h3 : 2'h0;
  assign T5702 = T5699[6'h2c:6'h2c];
  assign T5703 = $signed(T5704) / $signed(22'h100000);
  assign T5704 = $signed(31'h40c06355) * $signed(16'h0);
  assign twiddle4_3_359_imag = T5710 + T5705;
  assign T5705 = {T5708, T5706};
  assign T5706 = $signed(T5707) / $signed(22'h100000);
  assign T5707 = $signed(29'h15a3a741) * $signed(16'hffff);
  assign T5708 = T5709 ? 2'h3 : 2'h0;
  assign T5709 = T5706[6'h2c:6'h2c];
  assign T5710 = $signed(T5711) / $signed(22'h100000);
  assign T5711 = $signed(31'h40d81d61) * $signed(16'h0);
  assign T5712 = T2943[1'h0:1'h0];
  assign T5713 = T2943[1'h1:1'h1];
  assign T5714 = T2943[2'h2:2'h2];
  assign T5715 = T5784 ? T5750 : T5716;
  assign T5716 = T5749 ? T5733 : T5717;
  assign T5717 = T5732 ? twiddle4_3_361_imag : twiddle4_3_360_imag;
  assign twiddle4_3_360_imag = T5723 + T5718;
  assign T5718 = {T5721, T5719};
  assign T5719 = $signed(T5720) / $signed(22'h100000);
  assign T5720 = $signed(29'h150ef5de) * $signed(16'hffff);
  assign T5721 = T5722 ? 2'h3 : 2'h0;
  assign T5722 = T5719[6'h2c:6'h2c];
  assign T5723 = $signed(T5724) / $signed(22'h100000);
  assign T5724 = $signed(31'h40f1360c) * $signed(16'h0);
  assign twiddle4_3_361_imag = T5730 + T5725;
  assign T5725 = {T5728, T5726};
  assign T5726 = $signed(T5727) / $signed(22'h100000);
  assign T5727 = $signed(29'h147a813a) * $signed(16'hffff);
  assign T5728 = T5729 ? 2'h3 : 2'h0;
  assign T5729 = T5726[6'h2c:6'h2c];
  assign T5730 = $signed(T5731) / $signed(22'h100000);
  assign T5731 = $signed(31'h410bacc8) * $signed(16'h0);
  assign T5732 = T2943[1'h0:1'h0];
  assign T5733 = T5748 ? twiddle4_3_363_imag : twiddle4_3_362_imag;
  assign twiddle4_3_362_imag = T5739 + T5734;
  assign T5734 = {T5737, T5735};
  assign T5735 = $signed(T5736) / $signed(22'h100000);
  assign T5736 = $signed(29'h13e64c8c) * $signed(16'hffff);
  assign T5737 = T5738 ? 2'h3 : 2'h0;
  assign T5738 = T5735[6'h2c:6'h2c];
  assign T5739 = $signed(T5740) / $signed(22'h100000);
  assign T5740 = $signed(31'h41278105) * $signed(16'h0);
  assign twiddle4_3_363_imag = T5746 + T5741;
  assign T5741 = {T5744, T5742};
  assign T5742 = $signed(T5743) / $signed(22'h100000);
  assign T5743 = $signed(29'h13525b0c) * $signed(16'hffff);
  assign T5744 = T5745 ? 2'h3 : 2'h0;
  assign T5745 = T5742[6'h2c:6'h2c];
  assign T5746 = $signed(T5747) / $signed(22'h100000);
  assign T5747 = $signed(31'h4144b226) * $signed(16'h0);
  assign T5748 = T2943[1'h0:1'h0];
  assign T5749 = T2943[1'h1:1'h1];
  assign T5750 = T5783 ? T5767 : T5751;
  assign T5751 = T5766 ? twiddle4_3_365_imag : twiddle4_3_364_imag;
  assign twiddle4_3_364_imag = T5757 + T5752;
  assign T5752 = {T5755, T5753};
  assign T5753 = $signed(T5754) / $signed(22'h100000);
  assign T5754 = $signed(29'h12beafee) * $signed(16'hffff);
  assign T5755 = T5756 ? 2'h3 : 2'h0;
  assign T5756 = T5753[6'h2c:6'h2c];
  assign T5757 = $signed(T5758) / $signed(22'h100000);
  assign T5758 = $signed(31'h41633f8a) * $signed(16'h0);
  assign twiddle4_3_365_imag = T5764 + T5759;
  assign T5759 = {T5762, T5760};
  assign T5760 = $signed(T5761) / $signed(22'h100000);
  assign T5761 = $signed(29'h122b4e66) * $signed(16'hffff);
  assign T5762 = T5763 ? 2'h3 : 2'h0;
  assign T5763 = T5760[6'h2c:6'h2c];
  assign T5764 = $signed(T5765) / $signed(22'h100000);
  assign T5765 = $signed(31'h41832888) * $signed(16'h0);
  assign T5766 = T2943[1'h0:1'h0];
  assign T5767 = T5782 ? twiddle4_3_367_imag : twiddle4_3_366_imag;
  assign twiddle4_3_366_imag = T5773 + T5768;
  assign T5768 = {T5771, T5769};
  assign T5769 = $signed(T5770) / $signed(22'h100000);
  assign T5770 = $signed(29'h119839a7) * $signed(16'hffff);
  assign T5771 = T5772 ? 2'h3 : 2'h0;
  assign T5772 = T5769[6'h2c:6'h2c];
  assign T5773 = $signed(T5774) / $signed(22'h100000);
  assign T5774 = $signed(31'h41a46c6e) * $signed(16'h0);
  assign twiddle4_3_367_imag = T5780 + T5775;
  assign T5775 = {T5778, T5776};
  assign T5776 = $signed(T5777) / $signed(22'h100000);
  assign T5777 = $signed(29'h110574e1) * $signed(16'hffff);
  assign T5778 = T5779 ? 2'h3 : 2'h0;
  assign T5779 = T5776[6'h2c:6'h2c];
  assign T5780 = $signed(T5781) / $signed(22'h100000);
  assign T5781 = $signed(31'h41c70a84) * $signed(16'h0);
  assign T5782 = T2943[1'h0:1'h0];
  assign T5783 = T2943[1'h1:1'h1];
  assign T5784 = T2943[2'h2:2'h2];
  assign T5785 = T2943[2'h3:2'h3];
  assign T5786 = T5912 ? T5850 : T5787;
  assign T5787 = T5849 ? T5819 : T5788;
  assign T5788 = T5818 ? T5804 : T5789;
  assign T5789 = T5803 ? twiddle4_3_369_imag : twiddle4_3_368_imag;
  assign twiddle4_3_368_imag = T5795 + T5790;
  assign T5790 = {T5793, T5791};
  assign T5791 = $signed(T5792) / $signed(22'h100000);
  assign T5792 = $signed(29'h10730343) * $signed(16'hffff);
  assign T5793 = T5794 ? 2'h3 : 2'h0;
  assign T5794 = T5791[6'h2c:6'h2c];
  assign T5795 = $signed(T5796) / $signed(22'h100000);
  assign T5796 = $signed(31'h41eb0209) * $signed(16'h0);
  assign twiddle4_3_369_imag = T5801 + T5797;
  assign T5797 = {T5800, T5798};
  assign T5798 = $signed(T5799) / $signed(22'h100000);
  assign T5799 = $signed(30'h2fe0e7fa) * $signed(16'hffff);
  assign T5800 = T5798[6'h2d:6'h2d];
  assign T5801 = $signed(T5802) / $signed(22'h100000);
  assign T5802 = $signed(31'h42105236) * $signed(16'h0);
  assign T5803 = T2943[1'h0:1'h0];
  assign T5804 = T5817 ? twiddle4_3_371_imag : twiddle4_3_370_imag;
  assign twiddle4_3_370_imag = T5809 + T5805;
  assign T5805 = {T5808, T5806};
  assign T5806 = $signed(T5807) / $signed(22'h100000);
  assign T5807 = $signed(30'h2f4f2631) * $signed(16'hffff);
  assign T5808 = T5806[6'h2d:6'h2d];
  assign T5809 = $signed(T5810) / $signed(22'h100000);
  assign T5810 = $signed(31'h4236fa3c) * $signed(16'h0);
  assign twiddle4_3_371_imag = T5815 + T5811;
  assign T5811 = {T5814, T5812};
  assign T5812 = $signed(T5813) / $signed(22'h100000);
  assign T5813 = $signed(30'h2ebdc111) * $signed(16'hffff);
  assign T5814 = T5812[6'h2d:6'h2d];
  assign T5815 = $signed(T5816) / $signed(22'h100000);
  assign T5816 = $signed(31'h425ef943) * $signed(16'h0);
  assign T5817 = T2943[1'h0:1'h0];
  assign T5818 = T2943[1'h1:1'h1];
  assign T5819 = T5848 ? T5834 : T5820;
  assign T5820 = T5833 ? twiddle4_3_373_imag : twiddle4_3_372_imag;
  assign twiddle4_3_372_imag = T5825 + T5821;
  assign T5821 = {T5824, T5822};
  assign T5822 = $signed(T5823) / $signed(22'h100000);
  assign T5823 = $signed(30'h2e2cbbc1) * $signed(16'hffff);
  assign T5824 = T5822[6'h2d:6'h2d];
  assign T5825 = $signed(T5826) / $signed(22'h100000);
  assign T5826 = $signed(31'h42884e6f) * $signed(16'h0);
  assign twiddle4_3_373_imag = T5831 + T5827;
  assign T5827 = {T5830, T5828};
  assign T5828 = $signed(T5829) / $signed(22'h100000);
  assign T5829 = $signed(30'h2d9c1967) * $signed(16'hffff);
  assign T5830 = T5828[6'h2d:6'h2d];
  assign T5831 = $signed(T5832) / $signed(22'h100000);
  assign T5832 = $signed(31'h42b2f8d9) * $signed(16'h0);
  assign T5833 = T2943[1'h0:1'h0];
  assign T5834 = T5847 ? twiddle4_3_375_imag : twiddle4_3_374_imag;
  assign twiddle4_3_374_imag = T5839 + T5835;
  assign T5835 = {T5838, T5836};
  assign T5836 = $signed(T5837) / $signed(22'h100000);
  assign T5837 = $signed(30'h2d0bdd26) * $signed(16'hffff);
  assign T5838 = T5836[6'h2d:6'h2d];
  assign T5839 = $signed(T5840) / $signed(22'h100000);
  assign T5840 = $signed(31'h42def794) * $signed(16'h0);
  assign twiddle4_3_375_imag = T5845 + T5841;
  assign T5841 = {T5844, T5842};
  assign T5842 = $signed(T5843) / $signed(22'h100000);
  assign T5843 = $signed(30'h2c7c0a1d) * $signed(16'hffff);
  assign T5844 = T5842[6'h2d:6'h2d];
  assign T5845 = $signed(T5846) / $signed(22'h100000);
  assign T5846 = $signed(31'h430c49ad) * $signed(16'h0);
  assign T5847 = T2943[1'h0:1'h0];
  assign T5848 = T2943[1'h1:1'h1];
  assign T5849 = T2943[2'h2:2'h2];
  assign T5850 = T5911 ? T5881 : T5851;
  assign T5851 = T5880 ? T5866 : T5852;
  assign T5852 = T5865 ? twiddle4_3_377_imag : twiddle4_3_376_imag;
  assign twiddle4_3_376_imag = T5857 + T5853;
  assign T5853 = {T5856, T5854};
  assign T5854 = $signed(T5855) / $signed(22'h100000);
  assign T5855 = $signed(30'h2beca36c) * $signed(16'hffff);
  assign T5856 = T5854[6'h2d:6'h2d];
  assign T5857 = $signed(T5858) / $signed(22'h100000);
  assign T5858 = $signed(31'h433aee28) * $signed(16'h0);
  assign twiddle4_3_377_imag = T5863 + T5859;
  assign T5859 = {T5862, T5860};
  assign T5860 = $signed(T5861) / $signed(22'h100000);
  assign T5861 = $signed(30'h2b5dac2f) * $signed(16'hffff);
  assign T5862 = T5860[6'h2d:6'h2d];
  assign T5863 = $signed(T5864) / $signed(22'h100000);
  assign T5864 = $signed(31'h436ae401) * $signed(16'h0);
  assign T5865 = T2943[1'h0:1'h0];
  assign T5866 = T5879 ? twiddle4_3_379_imag : twiddle4_3_378_imag;
  assign twiddle4_3_378_imag = T5871 + T5867;
  assign T5867 = {T5870, T5868};
  assign T5868 = $signed(T5869) / $signed(22'h100000);
  assign T5869 = $signed(30'h2acf2780) * $signed(16'hffff);
  assign T5870 = T5868[6'h2d:6'h2d];
  assign T5871 = $signed(T5872) / $signed(22'h100000);
  assign T5872 = $signed(31'h439c2a30) * $signed(16'h0);
  assign twiddle4_3_379_imag = T5877 + T5873;
  assign T5873 = {T5876, T5874};
  assign T5874 = $signed(T5875) / $signed(22'h100000);
  assign T5875 = $signed(30'h2a411875) * $signed(16'hffff);
  assign T5876 = T5874[6'h2d:6'h2d];
  assign T5877 = $signed(T5878) / $signed(22'h100000);
  assign T5878 = $signed(31'h43cebfa1) * $signed(16'h0);
  assign T5879 = T2943[1'h0:1'h0];
  assign T5880 = T2943[1'h1:1'h1];
  assign T5881 = T5910 ? T5896 : T5882;
  assign T5882 = T5895 ? twiddle4_3_381_imag : twiddle4_3_380_imag;
  assign twiddle4_3_380_imag = T5887 + T5883;
  assign T5883 = {T5886, T5884};
  assign T5884 = $signed(T5885) / $signed(22'h100000);
  assign T5885 = $signed(30'h29b38223) * $signed(16'hffff);
  assign T5886 = T5884[6'h2d:6'h2d];
  assign T5887 = $signed(T5888) / $signed(22'h100000);
  assign T5888 = $signed(31'h4402a33c) * $signed(16'h0);
  assign twiddle4_3_381_imag = T5893 + T5889;
  assign T5889 = {T5892, T5890};
  assign T5890 = $signed(T5891) / $signed(22'h100000);
  assign T5891 = $signed(30'h2926679d) * $signed(16'hffff);
  assign T5892 = T5890[6'h2d:6'h2d];
  assign T5893 = $signed(T5894) / $signed(22'h100000);
  assign T5894 = $signed(31'h4437d3e2) * $signed(16'h0);
  assign T5895 = T2943[1'h0:1'h0];
  assign T5896 = T5909 ? twiddle4_3_383_imag : twiddle4_3_382_imag;
  assign twiddle4_3_382_imag = T5901 + T5897;
  assign T5897 = {T5900, T5898};
  assign T5898 = $signed(T5899) / $signed(22'h100000);
  assign T5899 = $signed(30'h2899cbf1) * $signed(16'hffff);
  assign T5900 = T5898[6'h2d:6'h2d];
  assign T5901 = $signed(T5902) / $signed(22'h100000);
  assign T5902 = $signed(31'h446e506a) * $signed(16'h0);
  assign twiddle4_3_383_imag = T5907 + T5903;
  assign T5903 = {T5906, T5904};
  assign T5904 = $signed(T5905) / $signed(22'h100000);
  assign T5905 = $signed(30'h280db22d) * $signed(16'hffff);
  assign T5906 = T5904[6'h2d:6'h2d];
  assign T5907 = $signed(T5908) / $signed(22'h100000);
  assign T5908 = $signed(31'h44a617a7) * $signed(16'h0);
  assign T5909 = T2943[1'h0:1'h0];
  assign T5910 = T2943[1'h1:1'h1];
  assign T5911 = T2943[2'h2:2'h2];
  assign T5912 = T2943[2'h3:2'h3];
  assign T5913 = T2943[3'h4:3'h4];
  assign T5914 = T2943[3'h5:3'h5];
  assign T5915 = T2943[3'h6:3'h6];
  assign T5916 = T6850 ? T6329 : T5917;
  assign T5917 = T6328 ? T6138 : T5918;
  assign T5918 = T6137 ? T6043 : T5919;
  assign T5919 = T6042 ? T5982 : T5920;
  assign T5920 = T5981 ? T5951 : T5921;
  assign T5921 = T5950 ? T5936 : T5922;
  assign T5922 = T5935 ? twiddle4_3_385_imag : twiddle4_3_384_imag;
  assign twiddle4_3_384_imag = T5927 + T5923;
  assign T5923 = {T5926, T5924};
  assign T5924 = $signed(T5925) / $signed(22'h100000);
  assign T5925 = $signed(30'h27821d5a) * $signed(16'hffff);
  assign T5926 = T5924[6'h2d:6'h2d];
  assign T5927 = $signed(T5928) / $signed(22'h100000);
  assign T5928 = $signed(31'h44df2862) * $signed(16'h0);
  assign twiddle4_3_385_imag = T5933 + T5929;
  assign T5929 = {T5932, T5930};
  assign T5930 = $signed(T5931) / $signed(22'h100000);
  assign T5931 = $signed(30'h26f7107f) * $signed(16'hffff);
  assign T5932 = T5930[6'h2d:6'h2d];
  assign T5933 = $signed(T5934) / $signed(22'h100000);
  assign T5934 = $signed(31'h4519815f) * $signed(16'h0);
  assign T5935 = T2943[1'h0:1'h0];
  assign T5936 = T5949 ? twiddle4_3_387_imag : twiddle4_3_386_imag;
  assign twiddle4_3_386_imag = T5941 + T5937;
  assign T5937 = {T5940, T5938};
  assign T5938 = $signed(T5939) / $signed(22'h100000);
  assign T5939 = $signed(30'h266c8e9f) * $signed(16'hffff);
  assign T5940 = T5938[6'h2d:6'h2d];
  assign T5941 = $signed(T5942) / $signed(22'h100000);
  assign T5942 = $signed(31'h4555215b) * $signed(16'h0);
  assign twiddle4_3_387_imag = T5947 + T5943;
  assign T5943 = {T5946, T5944};
  assign T5944 = $signed(T5945) / $signed(22'h100000);
  assign T5945 = $signed(30'h25e29abd) * $signed(16'hffff);
  assign T5946 = T5944[6'h2d:6'h2d];
  assign T5947 = $signed(T5948) / $signed(22'h100000);
  assign T5948 = $signed(31'h45920709) * $signed(16'h0);
  assign T5949 = T2943[1'h0:1'h0];
  assign T5950 = T2943[1'h1:1'h1];
  assign T5951 = T5980 ? T5966 : T5952;
  assign T5952 = T5965 ? twiddle4_3_389_imag : twiddle4_3_388_imag;
  assign twiddle4_3_388_imag = T5957 + T5953;
  assign T5953 = {T5956, T5954};
  assign T5954 = $signed(T5955) / $signed(22'h100000);
  assign T5955 = $signed(30'h255937d5) * $signed(16'hffff);
  assign T5956 = T5954[6'h2d:6'h2d];
  assign T5957 = $signed(T5958) / $signed(22'h100000);
  assign T5958 = $signed(31'h45d03118) * $signed(16'h0);
  assign twiddle4_3_389_imag = T5963 + T5959;
  assign T5959 = {T5962, T5960};
  assign T5960 = $signed(T5961) / $signed(22'h100000);
  assign T5961 = $signed(30'h24d068e3) * $signed(16'hffff);
  assign T5962 = T5960[6'h2d:6'h2d];
  assign T5963 = $signed(T5964) / $signed(22'h100000);
  assign T5964 = $signed(31'h460f9e2f) * $signed(16'h0);
  assign T5965 = T2943[1'h0:1'h0];
  assign T5966 = T5979 ? twiddle4_3_391_imag : twiddle4_3_390_imag;
  assign twiddle4_3_390_imag = T5971 + T5967;
  assign T5967 = {T5970, T5968};
  assign T5968 = $signed(T5969) / $signed(22'h100000);
  assign T5969 = $signed(30'h244830dd) * $signed(16'hffff);
  assign T5970 = T5968[6'h2d:6'h2d];
  assign T5971 = $signed(T5972) / $signed(22'h100000);
  assign T5972 = $signed(31'h46504ced) * $signed(16'h0);
  assign twiddle4_3_391_imag = T5977 + T5973;
  assign T5973 = {T5976, T5974};
  assign T5974 = $signed(T5975) / $signed(22'h100000);
  assign T5975 = $signed(30'h23c092b9) * $signed(16'hffff);
  assign T5976 = T5974[6'h2d:6'h2d];
  assign T5977 = $signed(T5978) / $signed(22'h100000);
  assign T5978 = $signed(31'h46923bec) * $signed(16'h0);
  assign T5979 = T2943[1'h0:1'h0];
  assign T5980 = T2943[1'h1:1'h1];
  assign T5981 = T2943[2'h2:2'h2];
  assign T5982 = T6041 ? T6013 : T5983;
  assign T5983 = T6012 ? T5998 : T5984;
  assign T5984 = T5997 ? twiddle4_3_393_imag : twiddle4_3_392_imag;
  assign twiddle4_3_392_imag = T5989 + T5985;
  assign T5985 = {T5988, T5986};
  assign T5986 = $signed(T5987) / $signed(22'h100000);
  assign T5987 = $signed(30'h23399167) * $signed(16'hffff);
  assign T5988 = T5986[6'h2d:6'h2d];
  assign T5989 = $signed(T5990) / $signed(22'h100000);
  assign T5990 = $signed(31'h46d569be) * $signed(16'h0);
  assign twiddle4_3_393_imag = T5995 + T5991;
  assign T5991 = {T5994, T5992};
  assign T5992 = $signed(T5993) / $signed(22'h100000);
  assign T5993 = $signed(30'h22b32fd5) * $signed(16'hffff);
  assign T5994 = T5992[6'h2d:6'h2d];
  assign T5995 = $signed(T5996) / $signed(22'h100000);
  assign T5996 = $signed(31'h4719d4ed) * $signed(16'h0);
  assign T5997 = T2943[1'h0:1'h0];
  assign T5998 = T6011 ? twiddle4_3_395_imag : twiddle4_3_394_imag;
  assign twiddle4_3_394_imag = T6003 + T5999;
  assign T5999 = {T6002, T6000};
  assign T6000 = $signed(T6001) / $signed(22'h100000);
  assign T6001 = $signed(30'h222d70ec) * $signed(16'hffff);
  assign T6002 = T6000[6'h2d:6'h2d];
  assign T6003 = $signed(T6004) / $signed(22'h100000);
  assign T6004 = $signed(31'h475f7bfe) * $signed(16'h0);
  assign twiddle4_3_395_imag = T6009 + T6005;
  assign T6005 = {T6008, T6006};
  assign T6006 = $signed(T6007) / $signed(22'h100000);
  assign T6007 = $signed(30'h21a85793) * $signed(16'hffff);
  assign T6008 = T6006[6'h2d:6'h2d];
  assign T6009 = $signed(T6010) / $signed(22'h100000);
  assign T6010 = $signed(31'h47a65d6e) * $signed(16'h0);
  assign T6011 = T2943[1'h0:1'h0];
  assign T6012 = T2943[1'h1:1'h1];
  assign T6013 = T6040 ? T6028 : T6014;
  assign T6014 = T6027 ? twiddle4_3_397_imag : twiddle4_3_396_imag;
  assign twiddle4_3_396_imag = T6019 + T6015;
  assign T6015 = {T6018, T6016};
  assign T6016 = $signed(T6017) / $signed(22'h100000);
  assign T6017 = $signed(30'h2123e6ae) * $signed(16'hffff);
  assign T6018 = T6016[6'h2d:6'h2d];
  assign T6019 = $signed(T6020) / $signed(22'h100000);
  assign T6020 = $signed(31'h47ee77b4) * $signed(16'h0);
  assign twiddle4_3_397_imag = T6025 + T6021;
  assign T6021 = {T6024, T6022};
  assign T6022 = $signed(T6023) / $signed(22'h100000);
  assign T6023 = $signed(30'h20a0211a) * $signed(16'hffff);
  assign T6024 = T6022[6'h2d:6'h2d];
  assign T6025 = $signed(T6026) / $signed(22'h100000);
  assign T6026 = $signed(31'h4837c93e) * $signed(16'h0);
  assign T6027 = T2943[1'h0:1'h0];
  assign T6028 = T6039 ? twiddle4_3_399_imag : twiddle4_3_398_imag;
  assign twiddle4_3_398_imag = T6033 + T6029;
  assign T6029 = {T6032, T6030};
  assign T6030 = $signed(T6031) / $signed(22'h100000);
  assign T6031 = $signed(30'h201d09b5) * $signed(16'hffff);
  assign T6032 = T6030[6'h2d:6'h2d];
  assign T6033 = $signed(T6034) / $signed(22'h100000);
  assign T6034 = $signed(31'h48825077) * $signed(16'h0);
  assign twiddle4_3_399_imag = T6037 + T6035;
  assign T6035 = $signed(T6036) / $signed(22'h100000);
  assign T6036 = $signed(31'h5f9aa355) * $signed(16'hffff);
  assign T6037 = $signed(T6038) / $signed(22'h100000);
  assign T6038 = $signed(31'h48ce0bc1) * $signed(16'h0);
  assign T6039 = T2943[1'h0:1'h0];
  assign T6040 = T2943[1'h1:1'h1];
  assign T6041 = T2943[2'h2:2'h2];
  assign T6042 = T2943[2'h3:2'h3];
  assign T6043 = T6136 ? T6090 : T6044;
  assign T6044 = T6089 ? T6067 : T6045;
  assign T6045 = T6066 ? T6056 : T6046;
  assign T6046 = T6055 ? twiddle4_3_401_imag : twiddle4_3_400_imag;
  assign twiddle4_3_400_imag = T6049 + T6047;
  assign T6047 = $signed(T6048) / $signed(22'h100000);
  assign T6048 = $signed(31'h5f18f0ce) * $signed(16'hffff);
  assign T6049 = $signed(T6050) / $signed(22'h100000);
  assign T6050 = $signed(31'h491af976) * $signed(16'h0);
  assign twiddle4_3_401_imag = T6053 + T6051;
  assign T6051 = $signed(T6052) / $signed(22'h100000);
  assign T6052 = $signed(31'h5e97f4f1) * $signed(16'hffff);
  assign T6053 = $signed(T6054) / $signed(22'h100000);
  assign T6054 = $signed(31'h496917ed) * $signed(16'h0);
  assign T6055 = T2943[1'h0:1'h0];
  assign T6056 = T6065 ? twiddle4_3_403_imag : twiddle4_3_402_imag;
  assign twiddle4_3_402_imag = T6059 + T6057;
  assign T6057 = $signed(T6058) / $signed(22'h100000);
  assign T6058 = $signed(31'h5e17b28a) * $signed(16'hffff);
  assign T6059 = $signed(T6060) / $signed(22'h100000);
  assign T6060 = $signed(31'h49b86572) * $signed(16'h0);
  assign twiddle4_3_403_imag = T6063 + T6061;
  assign T6061 = $signed(T6062) / $signed(22'h100000);
  assign T6062 = $signed(31'h5d982c61) * $signed(16'hffff);
  assign T6063 = $signed(T6064) / $signed(22'h100000);
  assign T6064 = $signed(31'h4a08e04f) * $signed(16'h0);
  assign T6065 = T2943[1'h0:1'h0];
  assign T6066 = T2943[1'h1:1'h1];
  assign T6067 = T6088 ? T6078 : T6068;
  assign T6068 = T6077 ? twiddle4_3_405_imag : twiddle4_3_404_imag;
  assign twiddle4_3_404_imag = T6071 + T6069;
  assign T6069 = $signed(T6070) / $signed(22'h100000);
  assign T6070 = $signed(31'h5d196539) * $signed(16'hffff);
  assign T6071 = $signed(T6072) / $signed(22'h100000);
  assign T6072 = $signed(31'h4a5a86c4) * $signed(16'h0);
  assign twiddle4_3_405_imag = T6075 + T6073;
  assign T6073 = $signed(T6074) / $signed(22'h100000);
  assign T6074 = $signed(31'h5c9b5fd2) * $signed(16'hffff);
  assign T6075 = $signed(T6076) / $signed(22'h100000);
  assign T6076 = $signed(31'h4aad570c) * $signed(16'h0);
  assign T6077 = T2943[1'h0:1'h0];
  assign T6078 = T6087 ? twiddle4_3_407_imag : twiddle4_3_406_imag;
  assign twiddle4_3_406_imag = T6081 + T6079;
  assign T6079 = $signed(T6080) / $signed(22'h100000);
  assign T6080 = $signed(31'h5c1e1ee9) * $signed(16'hffff);
  assign T6081 = $signed(T6082) / $signed(22'h100000);
  assign T6082 = $signed(31'h4b014f5b) * $signed(16'h0);
  assign twiddle4_3_407_imag = T6085 + T6083;
  assign T6083 = $signed(T6084) / $signed(22'h100000);
  assign T6084 = $signed(31'h5ba1a534) * $signed(16'hffff);
  assign T6085 = $signed(T6086) / $signed(22'h100000);
  assign T6086 = $signed(31'h4b566ddf) * $signed(16'h0);
  assign T6087 = T2943[1'h0:1'h0];
  assign T6088 = T2943[1'h1:1'h1];
  assign T6089 = T2943[2'h2:2'h2];
  assign T6090 = T6135 ? T6113 : T6091;
  assign T6091 = T6112 ? T6102 : T6092;
  assign T6092 = T6101 ? twiddle4_3_409_imag : twiddle4_3_408_imag;
  assign twiddle4_3_408_imag = T6095 + T6093;
  assign T6093 = $signed(T6094) / $signed(22'h100000);
  assign T6094 = $signed(31'h5b25f567) * $signed(16'hffff);
  assign T6095 = $signed(T6096) / $signed(22'h100000);
  assign T6096 = $signed(31'h4bacb0c0) * $signed(16'h0);
  assign twiddle4_3_409_imag = T6099 + T6097;
  assign T6097 = $signed(T6098) / $signed(22'h100000);
  assign T6098 = $signed(31'h5aab1230) * $signed(16'hffff);
  assign T6099 = $signed(T6100) / $signed(22'h100000);
  assign T6100 = $signed(31'h4c04161e) * $signed(16'h0);
  assign T6101 = T2943[1'h0:1'h0];
  assign T6102 = T6111 ? twiddle4_3_411_imag : twiddle4_3_410_imag;
  assign twiddle4_3_410_imag = T6105 + T6103;
  assign T6103 = $signed(T6104) / $signed(22'h100000);
  assign T6104 = $signed(31'h5a30fe39) * $signed(16'hffff);
  assign T6105 = $signed(T6106) / $signed(22'h100000);
  assign T6106 = $signed(31'h4c5c9c15) * $signed(16'h0);
  assign twiddle4_3_411_imag = T6109 + T6107;
  assign T6107 = $signed(T6108) / $signed(22'h100000);
  assign T6108 = $signed(31'h59b7bc28) * $signed(16'hffff);
  assign T6109 = $signed(T6110) / $signed(22'h100000);
  assign T6110 = $signed(31'h4cb640b8) * $signed(16'h0);
  assign T6111 = T2943[1'h0:1'h0];
  assign T6112 = T2943[1'h1:1'h1];
  assign T6113 = T6134 ? T6124 : T6114;
  assign T6114 = T6123 ? twiddle4_3_413_imag : twiddle4_3_412_imag;
  assign twiddle4_3_412_imag = T6117 + T6115;
  assign T6115 = $signed(T6116) / $signed(22'h100000);
  assign T6116 = $signed(31'h593f4e9e) * $signed(16'hffff);
  assign T6117 = $signed(T6118) / $signed(22'h100000);
  assign T6118 = $signed(31'h4d110217) * $signed(16'h0);
  assign twiddle4_3_413_imag = T6121 + T6119;
  assign T6119 = $signed(T6120) / $signed(22'h100000);
  assign T6120 = $signed(31'h58c7b839) * $signed(16'hffff);
  assign T6121 = $signed(T6122) / $signed(22'h100000);
  assign T6122 = $signed(31'h4d6cde39) * $signed(16'h0);
  assign T6123 = T2943[1'h0:1'h0];
  assign T6124 = T6133 ? twiddle4_3_415_imag : twiddle4_3_414_imag;
  assign twiddle4_3_414_imag = T6127 + T6125;
  assign T6125 = $signed(T6126) / $signed(22'h100000);
  assign T6126 = $signed(31'h5850fb8f) * $signed(16'hffff);
  assign T6127 = $signed(T6128) / $signed(22'h100000);
  assign T6128 = $signed(31'h4dc9d321) * $signed(16'h0);
  assign twiddle4_3_415_imag = T6131 + T6129;
  assign T6129 = $signed(T6130) / $signed(22'h100000);
  assign T6130 = $signed(31'h57db1b34) * $signed(16'hffff);
  assign T6131 = $signed(T6132) / $signed(22'h100000);
  assign T6132 = $signed(31'h4e27deca) * $signed(16'h0);
  assign T6133 = T2943[1'h0:1'h0];
  assign T6134 = T2943[1'h1:1'h1];
  assign T6135 = T2943[2'h2:2'h2];
  assign T6136 = T2943[2'h3:2'h3];
  assign T6137 = T2943[3'h4:3'h4];
  assign T6138 = T6327 ? T6233 : T6139;
  assign T6139 = T6232 ? T6186 : T6140;
  assign T6140 = T6185 ? T6163 : T6141;
  assign T6141 = T6162 ? T6152 : T6142;
  assign T6142 = T6151 ? twiddle4_3_417_imag : twiddle4_3_416_imag;
  assign twiddle4_3_416_imag = T6145 + T6143;
  assign T6143 = $signed(T6144) / $signed(22'h100000);
  assign T6144 = $signed(31'h576619b6) * $signed(16'hffff);
  assign T6145 = $signed(T6146) / $signed(22'h100000);
  assign T6146 = $signed(31'h4e86ff2a) * $signed(16'h0);
  assign twiddle4_3_417_imag = T6149 + T6147;
  assign T6147 = $signed(T6148) / $signed(22'h100000);
  assign T6148 = $signed(31'h56f1f9a0) * $signed(16'hffff);
  assign T6149 = $signed(T6150) / $signed(22'h100000);
  assign T6150 = $signed(31'h4ee73232) * $signed(16'h0);
  assign T6151 = T2943[1'h0:1'h0];
  assign T6152 = T6161 ? twiddle4_3_419_imag : twiddle4_3_418_imag;
  assign twiddle4_3_418_imag = T6155 + T6153;
  assign T6153 = $signed(T6154) / $signed(22'h100000);
  assign T6154 = $signed(31'h567ebd75) * $signed(16'hffff);
  assign T6155 = $signed(T6156) / $signed(22'h100000);
  assign T6156 = $signed(31'h4f4875cb) * $signed(16'h0);
  assign twiddle4_3_419_imag = T6159 + T6157;
  assign T6157 = $signed(T6158) / $signed(22'h100000);
  assign T6158 = $signed(31'h560c67b5) * $signed(16'hffff);
  assign T6159 = $signed(T6160) / $signed(22'h100000);
  assign T6160 = $signed(31'h4faac7d9) * $signed(16'h0);
  assign T6161 = T2943[1'h0:1'h0];
  assign T6162 = T2943[1'h1:1'h1];
  assign T6163 = T6184 ? T6174 : T6164;
  assign T6164 = T6173 ? twiddle4_3_421_imag : twiddle4_3_420_imag;
  assign twiddle4_3_420_imag = T6167 + T6165;
  assign T6165 = $signed(T6166) / $signed(22'h100000);
  assign T6166 = $signed(31'h559afadb) * $signed(16'hffff);
  assign T6167 = $signed(T6168) / $signed(22'h100000);
  assign T6168 = $signed(31'h500e263a) * $signed(16'h0);
  assign twiddle4_3_421_imag = T6171 + T6169;
  assign T6169 = $signed(T6170) / $signed(22'h100000);
  assign T6170 = $signed(31'h552a795d) * $signed(16'hffff);
  assign T6171 = $signed(T6172) / $signed(22'h100000);
  assign T6172 = $signed(31'h50728ec7) * $signed(16'h0);
  assign T6173 = T2943[1'h0:1'h0];
  assign T6174 = T6183 ? twiddle4_3_423_imag : twiddle4_3_422_imag;
  assign twiddle4_3_422_imag = T6177 + T6175;
  assign T6175 = $signed(T6176) / $signed(22'h100000);
  assign T6176 = $signed(31'h54bae5ac) * $signed(16'hffff);
  assign T6177 = $signed(T6178) / $signed(22'h100000);
  assign T6178 = $signed(31'h50d7ff52) * $signed(16'h0);
  assign twiddle4_3_423_imag = T6181 + T6179;
  assign T6179 = $signed(T6180) / $signed(22'h100000);
  assign T6180 = $signed(31'h544c4232) * $signed(16'hffff);
  assign T6181 = $signed(T6182) / $signed(22'h100000);
  assign T6182 = $signed(31'h513e75a8) * $signed(16'h0);
  assign T6183 = T2943[1'h0:1'h0];
  assign T6184 = T2943[1'h1:1'h1];
  assign T6185 = T2943[2'h2:2'h2];
  assign T6186 = T6231 ? T6209 : T6187;
  assign T6187 = T6208 ? T6198 : T6188;
  assign T6188 = T6197 ? twiddle4_3_425_imag : twiddle4_3_424_imag;
  assign twiddle4_3_424_imag = T6191 + T6189;
  assign T6189 = $signed(T6190) / $signed(22'h100000);
  assign T6190 = $signed(31'h53de9156) * $signed(16'hffff);
  assign T6191 = $signed(T6192) / $signed(22'h100000);
  assign T6192 = $signed(31'h51a5ef91) * $signed(16'h0);
  assign twiddle4_3_425_imag = T6195 + T6193;
  assign T6193 = $signed(T6194) / $signed(22'h100000);
  assign T6194 = $signed(31'h5371d57a) * $signed(16'hffff);
  assign T6195 = $signed(T6196) / $signed(22'h100000);
  assign T6196 = $signed(31'h520e6acd) * $signed(16'h0);
  assign T6197 = T2943[1'h0:1'h0];
  assign T6198 = T6207 ? twiddle4_3_427_imag : twiddle4_3_426_imag;
  assign twiddle4_3_426_imag = T6201 + T6199;
  assign T6199 = $signed(T6200) / $signed(22'h100000);
  assign T6200 = $signed(31'h530610f7) * $signed(16'hffff);
  assign T6201 = $signed(T6202) / $signed(22'h100000);
  assign T6202 = $signed(31'h5277e519) * $signed(16'h0);
  assign twiddle4_3_427_imag = T6205 + T6203;
  assign T6203 = $signed(T6204) / $signed(22'h100000);
  assign T6204 = $signed(31'h529b4626) * $signed(16'hffff);
  assign T6205 = $signed(T6206) / $signed(22'h100000);
  assign T6206 = $signed(31'h52e25c2b) * $signed(16'h0);
  assign T6207 = T2943[1'h0:1'h0];
  assign T6208 = T2943[1'h1:1'h1];
  assign T6209 = T6230 ? T6220 : T6210;
  assign T6210 = T6219 ? twiddle4_3_429_imag : twiddle4_3_428_imag;
  assign twiddle4_3_428_imag = T6213 + T6211;
  assign T6211 = $signed(T6212) / $signed(22'h100000);
  assign T6212 = $signed(31'h52317757) * $signed(16'hffff);
  assign T6213 = $signed(T6214) / $signed(22'h100000);
  assign T6214 = $signed(31'h534dcdb5) * $signed(16'h0);
  assign twiddle4_3_429_imag = T6217 + T6215;
  assign T6215 = $signed(T6216) / $signed(22'h100000);
  assign T6216 = $signed(31'h51c8a6d4) * $signed(16'hffff);
  assign T6217 = $signed(T6218) / $signed(22'h100000);
  assign T6218 = $signed(31'h53ba3761) * $signed(16'h0);
  assign T6219 = T2943[1'h0:1'h0];
  assign T6220 = T6229 ? twiddle4_3_431_imag : twiddle4_3_430_imag;
  assign twiddle4_3_430_imag = T6223 + T6221;
  assign T6221 = $signed(T6222) / $signed(22'h100000);
  assign T6222 = $signed(31'h5160d6e5) * $signed(16'hffff);
  assign T6223 = $signed(T6224) / $signed(22'h100000);
  assign T6224 = $signed(31'h542796d5) * $signed(16'h0);
  assign twiddle4_3_431_imag = T6227 + T6225;
  assign T6225 = $signed(T6226) / $signed(22'h100000);
  assign T6226 = $signed(31'h50fa09c9) * $signed(16'hffff);
  assign T6227 = $signed(T6228) / $signed(22'h100000);
  assign T6228 = $signed(31'h5495e9b4) * $signed(16'h0);
  assign T6229 = T2943[1'h0:1'h0];
  assign T6230 = T2943[1'h1:1'h1];
  assign T6231 = T2943[2'h2:2'h2];
  assign T6232 = T2943[2'h3:2'h3];
  assign T6233 = T6326 ? T6280 : T6234;
  assign T6234 = T6279 ? T6257 : T6235;
  assign T6235 = T6256 ? T6246 : T6236;
  assign T6236 = T6245 ? twiddle4_3_433_imag : twiddle4_3_432_imag;
  assign twiddle4_3_432_imag = T6239 + T6237;
  assign T6237 = $signed(T6238) / $signed(22'h100000);
  assign T6238 = $signed(31'h509441bc) * $signed(16'hffff);
  assign T6239 = $signed(T6240) / $signed(22'h100000);
  assign T6240 = $signed(31'h55052d97) * $signed(16'h0);
  assign twiddle4_3_433_imag = T6243 + T6241;
  assign T6241 = $signed(T6242) / $signed(22'h100000);
  assign T6242 = $signed(31'h502f80f1) * $signed(16'hffff);
  assign T6243 = $signed(T6244) / $signed(22'h100000);
  assign T6244 = $signed(31'h55756016) * $signed(16'h0);
  assign T6245 = T2943[1'h0:1'h0];
  assign T6246 = T6255 ? twiddle4_3_435_imag : twiddle4_3_434_imag;
  assign twiddle4_3_434_imag = T6249 + T6247;
  assign T6247 = $signed(T6248) / $signed(22'h100000);
  assign T6248 = $signed(31'h4fcbc999) * $signed(16'hffff);
  assign T6249 = $signed(T6250) / $signed(22'h100000);
  assign T6250 = $signed(31'h55e67ec2) * $signed(16'h0);
  assign twiddle4_3_435_imag = T6253 + T6251;
  assign T6251 = $signed(T6252) / $signed(22'h100000);
  assign T6252 = $signed(31'h4f691ddd) * $signed(16'hffff);
  assign T6253 = $signed(T6254) / $signed(22'h100000);
  assign T6254 = $signed(31'h56588726) * $signed(16'h0);
  assign T6255 = T2943[1'h0:1'h0];
  assign T6256 = T2943[1'h1:1'h1];
  assign T6257 = T6278 ? T6268 : T6258;
  assign T6258 = T6267 ? twiddle4_3_437_imag : twiddle4_3_436_imag;
  assign twiddle4_3_436_imag = T6261 + T6259;
  assign T6259 = $signed(T6260) / $signed(22'h100000);
  assign T6260 = $signed(31'h4f077fe1) * $signed(16'hffff);
  assign T6261 = $signed(T6262) / $signed(22'h100000);
  assign T6262 = $signed(31'h56cb76c9) * $signed(16'h0);
  assign twiddle4_3_437_imag = T6265 + T6263;
  assign T6263 = $signed(T6264) / $signed(22'h100000);
  assign T6264 = $signed(31'h4ea6f1c3) * $signed(16'hffff);
  assign T6265 = $signed(T6266) / $signed(22'h100000);
  assign T6266 = $signed(31'h573f4b2e) * $signed(16'h0);
  assign T6267 = T2943[1'h0:1'h0];
  assign T6268 = T6277 ? twiddle4_3_439_imag : twiddle4_3_438_imag;
  assign twiddle4_3_438_imag = T6271 + T6269;
  assign T6269 = $signed(T6270) / $signed(22'h100000);
  assign T6270 = $signed(31'h4e47759a) * $signed(16'hffff);
  assign T6271 = $signed(T6272) / $signed(22'h100000);
  assign T6272 = $signed(31'h57b401d1) * $signed(16'h0);
  assign twiddle4_3_439_imag = T6275 + T6273;
  assign T6273 = $signed(T6274) / $signed(22'h100000);
  assign T6274 = $signed(31'h4de90d7a) * $signed(16'hffff);
  assign T6275 = $signed(T6276) / $signed(22'h100000);
  assign T6276 = $signed(31'h5829982b) * $signed(16'h0);
  assign T6277 = T2943[1'h0:1'h0];
  assign T6278 = T2943[1'h1:1'h1];
  assign T6279 = T2943[2'h2:2'h2];
  assign T6280 = T6325 ? T6303 : T6281;
  assign T6281 = T6302 ? T6292 : T6282;
  assign T6282 = T6291 ? twiddle4_3_441_imag : twiddle4_3_440_imag;
  assign twiddle4_3_440_imag = T6285 + T6283;
  assign T6283 = $signed(T6284) / $signed(22'h100000);
  assign T6284 = $signed(31'h4d8bbb6d) * $signed(16'hffff);
  assign T6285 = $signed(T6286) / $signed(22'h100000);
  assign T6286 = $signed(31'h58a00bae) * $signed(16'h0);
  assign twiddle4_3_441_imag = T6289 + T6287;
  assign T6287 = $signed(T6288) / $signed(22'h100000);
  assign T6288 = $signed(31'h4d2f817b) * $signed(16'hffff);
  assign T6289 = $signed(T6290) / $signed(22'h100000);
  assign T6290 = $signed(31'h591759c9) * $signed(16'h0);
  assign T6291 = T2943[1'h0:1'h0];
  assign T6292 = T6301 ? twiddle4_3_443_imag : twiddle4_3_442_imag;
  assign twiddle4_3_442_imag = T6295 + T6293;
  assign T6293 = $signed(T6294) / $signed(22'h100000);
  assign T6294 = $signed(31'h4cd461a3) * $signed(16'hffff);
  assign T6295 = $signed(T6296) / $signed(22'h100000);
  assign T6296 = $signed(31'h598f7fe6) * $signed(16'h0);
  assign twiddle4_3_443_imag = T6299 + T6297;
  assign T6297 = $signed(T6298) / $signed(22'h100000);
  assign T6298 = $signed(31'h4c7a5ddf) * $signed(16'hffff);
  assign T6299 = $signed(T6300) / $signed(22'h100000);
  assign T6300 = $signed(31'h5a087b6a) * $signed(16'h0);
  assign T6301 = T2943[1'h0:1'h0];
  assign T6302 = T2943[1'h1:1'h1];
  assign T6303 = T6324 ? T6314 : T6304;
  assign T6304 = T6313 ? twiddle4_3_445_imag : twiddle4_3_444_imag;
  assign twiddle4_3_444_imag = T6307 + T6305;
  assign T6305 = $signed(T6306) / $signed(22'h100000);
  assign T6306 = $signed(31'h4c217822) * $signed(16'hffff);
  assign T6307 = $signed(T6308) / $signed(22'h100000);
  assign T6308 = $signed(31'h5a8249b5) * $signed(16'h0);
  assign twiddle4_3_445_imag = T6311 + T6309;
  assign T6309 = $signed(T6310) / $signed(22'h100000);
  assign T6310 = $signed(31'h4bc9b25b) * $signed(16'hffff);
  assign T6311 = $signed(T6312) / $signed(22'h100000);
  assign T6312 = $signed(31'h5afce822) * $signed(16'h0);
  assign T6313 = T2943[1'h0:1'h0];
  assign T6314 = T6323 ? twiddle4_3_447_imag : twiddle4_3_446_imag;
  assign twiddle4_3_446_imag = T6317 + T6315;
  assign T6315 = $signed(T6316) / $signed(22'h100000);
  assign T6316 = $signed(31'h4b730e70) * $signed(16'hffff);
  assign T6317 = $signed(T6318) / $signed(22'h100000);
  assign T6318 = $signed(31'h5b785409) * $signed(16'h0);
  assign twiddle4_3_447_imag = T6321 + T6319;
  assign T6319 = $signed(T6320) / $signed(22'h100000);
  assign T6320 = $signed(31'h4b1d8e43) * $signed(16'hffff);
  assign T6321 = $signed(T6322) / $signed(22'h100000);
  assign T6322 = $signed(31'h5bf48abe) * $signed(16'h0);
  assign T6323 = T2943[1'h0:1'h0];
  assign T6324 = T2943[1'h1:1'h1];
  assign T6325 = T2943[2'h2:2'h2];
  assign T6326 = T2943[2'h3:2'h3];
  assign T6327 = T2943[3'h4:3'h4];
  assign T6328 = T2943[3'h5:3'h5];
  assign T6329 = T6849 ? T6568 : T6330;
  assign T6330 = T6567 ? T6441 : T6331;
  assign T6331 = T6440 ? T6378 : T6332;
  assign T6332 = T6377 ? T6355 : T6333;
  assign T6333 = T6354 ? T6344 : T6334;
  assign T6334 = T6343 ? twiddle4_3_449_imag : twiddle4_3_448_imag;
  assign twiddle4_3_448_imag = T6337 + T6335;
  assign T6335 = $signed(T6336) / $signed(22'h100000);
  assign T6336 = $signed(31'h4ac933ae) * $signed(16'hffff);
  assign T6337 = $signed(T6338) / $signed(22'h100000);
  assign T6338 = $signed(31'h5c71898d) * $signed(16'h0);
  assign twiddle4_3_449_imag = T6341 + T6339;
  assign T6339 = $signed(T6340) / $signed(22'h100000);
  assign T6340 = $signed(31'h4a760086) * $signed(16'hffff);
  assign T6341 = $signed(T6342) / $signed(22'h100000);
  assign T6342 = $signed(31'h5cef4dc2) * $signed(16'h0);
  assign T6343 = T2943[1'h0:1'h0];
  assign T6344 = T6353 ? twiddle4_3_451_imag : twiddle4_3_450_imag;
  assign twiddle4_3_450_imag = T6347 + T6345;
  assign T6345 = $signed(T6346) / $signed(22'h100000);
  assign T6346 = $signed(31'h4a23f698) * $signed(16'hffff);
  assign T6347 = $signed(T6348) / $signed(22'h100000);
  assign T6348 = $signed(31'h5d6dd4a2) * $signed(16'h0);
  assign twiddle4_3_451_imag = T6351 + T6349;
  assign T6349 = $signed(T6350) / $signed(22'h100000);
  assign T6350 = $signed(31'h49d317ac) * $signed(16'hffff);
  assign T6351 = $signed(T6352) / $signed(22'h100000);
  assign T6352 = $signed(31'h5ded1b6f) * $signed(16'h0);
  assign T6353 = T2943[1'h0:1'h0];
  assign T6354 = T2943[1'h1:1'h1];
  assign T6355 = T6376 ? T6366 : T6356;
  assign T6356 = T6365 ? twiddle4_3_453_imag : twiddle4_3_452_imag;
  assign twiddle4_3_452_imag = T6359 + T6357;
  assign T6357 = $signed(T6358) / $signed(22'h100000);
  assign T6358 = $signed(31'h49836583) * $signed(16'hffff);
  assign T6359 = $signed(T6360) / $signed(22'h100000);
  assign T6360 = $signed(31'h5e6d1f66) * $signed(16'h0);
  assign twiddle4_3_453_imag = T6363 + T6361;
  assign T6361 = $signed(T6362) / $signed(22'h100000);
  assign T6362 = $signed(31'h4934e1d7) * $signed(16'hffff);
  assign T6363 = $signed(T6364) / $signed(22'h100000);
  assign T6364 = $signed(31'h5eedddc0) * $signed(16'h0);
  assign T6365 = T2943[1'h0:1'h0];
  assign T6366 = T6375 ? twiddle4_3_455_imag : twiddle4_3_454_imag;
  assign twiddle4_3_454_imag = T6369 + T6367;
  assign T6367 = $signed(T6368) / $signed(22'h100000);
  assign T6368 = $signed(31'h48e78e5c) * $signed(16'hffff);
  assign T6369 = $signed(T6370) / $signed(22'h100000);
  assign T6370 = $signed(31'h5f6f53b3) * $signed(16'h0);
  assign twiddle4_3_455_imag = T6373 + T6371;
  assign T6371 = $signed(T6372) / $signed(22'h100000);
  assign T6372 = $signed(31'h489b6cbf) * $signed(16'hffff);
  assign T6373 = $signed(T6374) / $signed(22'h100000);
  assign T6374 = $signed(31'h5ff17e70) * $signed(16'h0);
  assign T6375 = T2943[1'h0:1'h0];
  assign T6376 = T2943[1'h1:1'h1];
  assign T6377 = T2943[2'h2:2'h2];
  assign T6378 = T6439 ? T6409 : T6379;
  assign T6379 = T6408 ? T6394 : T6380;
  assign T6380 = T6393 ? twiddle4_3_457_imag : twiddle4_3_456_imag;
  assign twiddle4_3_456_imag = T6383 + T6381;
  assign T6381 = $signed(T6382) / $signed(22'h100000);
  assign T6382 = $signed(31'h48507ea8) * $signed(16'hffff);
  assign T6383 = {T6386, T6384};
  assign T6384 = $signed(T6385) / $signed(22'h100000);
  assign T6385 = $signed(30'h20745b25) * $signed(16'h0);
  assign T6386 = T6384[6'h2d:6'h2d];
  assign twiddle4_3_457_imag = T6389 + T6387;
  assign T6387 = $signed(T6388) / $signed(22'h100000);
  assign T6388 = $signed(31'h4806c5b5) * $signed(16'hffff);
  assign T6389 = {T6392, T6390};
  assign T6390 = $signed(T6391) / $signed(22'h100000);
  assign T6391 = $signed(30'h20f7e6fa) * $signed(16'h0);
  assign T6392 = T6390[6'h2d:6'h2d];
  assign T6393 = T2943[1'h0:1'h0];
  assign T6394 = T6407 ? twiddle4_3_459_imag : twiddle4_3_458_imag;
  assign twiddle4_3_458_imag = T6397 + T6395;
  assign T6395 = $signed(T6396) / $signed(22'h100000);
  assign T6396 = $signed(31'h47be4381) * $signed(16'hffff);
  assign T6397 = {T6400, T6398};
  assign T6398 = $signed(T6399) / $signed(22'h100000);
  assign T6399 = $signed(30'h217c1f16) * $signed(16'h0);
  assign T6400 = T6398[6'h2d:6'h2d];
  assign twiddle4_3_459_imag = T6403 + T6401;
  assign T6401 = $signed(T6402) / $signed(22'h100000);
  assign T6402 = $signed(31'h4776f99e) * $signed(16'hffff);
  assign T6403 = {T6406, T6404};
  assign T6404 = $signed(T6405) / $signed(22'h100000);
  assign T6405 = $signed(30'h2201009a) * $signed(16'h0);
  assign T6406 = T6404[6'h2d:6'h2d];
  assign T6407 = T2943[1'h0:1'h0];
  assign T6408 = T2943[1'h1:1'h1];
  assign T6409 = T6438 ? T6424 : T6410;
  assign T6410 = T6423 ? twiddle4_3_461_imag : twiddle4_3_460_imag;
  assign twiddle4_3_460_imag = T6413 + T6411;
  assign T6411 = $signed(T6412) / $signed(22'h100000);
  assign T6412 = $signed(31'h4730e997) * $signed(16'hffff);
  assign T6413 = {T6416, T6414};
  assign T6414 = $signed(T6415) / $signed(22'h100000);
  assign T6415 = $signed(30'h228688a5) * $signed(16'h0);
  assign T6416 = T6414[6'h2d:6'h2d];
  assign twiddle4_3_461_imag = T6419 + T6417;
  assign T6417 = $signed(T6418) / $signed(22'h100000);
  assign T6418 = $signed(31'h46ec14f2) * $signed(16'hffff);
  assign T6419 = {T6422, T6420};
  assign T6420 = $signed(T6421) / $signed(22'h100000);
  assign T6421 = $signed(30'h230cb452) * $signed(16'h0);
  assign T6422 = T6420[6'h2d:6'h2d];
  assign T6423 = T2943[1'h0:1'h0];
  assign T6424 = T6437 ? twiddle4_3_463_imag : twiddle4_3_462_imag;
  assign twiddle4_3_462_imag = T6427 + T6425;
  assign T6425 = $signed(T6426) / $signed(22'h100000);
  assign T6426 = $signed(31'h46a87d2d) * $signed(16'hffff);
  assign T6427 = {T6430, T6428};
  assign T6428 = $signed(T6429) / $signed(22'h100000);
  assign T6429 = $signed(30'h239380b7) * $signed(16'h0);
  assign T6430 = T6428[6'h2d:6'h2d];
  assign twiddle4_3_463_imag = T6433 + T6431;
  assign T6431 = $signed(T6432) / $signed(22'h100000);
  assign T6432 = $signed(31'h466623bf) * $signed(16'hffff);
  assign T6433 = {T6436, T6434};
  assign T6434 = $signed(T6435) / $signed(22'h100000);
  assign T6435 = $signed(30'h241aeae9) * $signed(16'h0);
  assign T6436 = T6434[6'h2d:6'h2d];
  assign T6437 = T2943[1'h0:1'h0];
  assign T6438 = T2943[1'h1:1'h1];
  assign T6439 = T2943[2'h2:2'h2];
  assign T6440 = T2943[2'h3:2'h3];
  assign T6441 = T6566 ? T6504 : T6442;
  assign T6442 = T6503 ? T6473 : T6443;
  assign T6443 = T6472 ? T6458 : T6444;
  assign T6444 = T6457 ? twiddle4_3_465_imag : twiddle4_3_464_imag;
  assign twiddle4_3_464_imag = T6447 + T6445;
  assign T6445 = $signed(T6446) / $signed(22'h100000);
  assign T6446 = $signed(31'h46250a18) * $signed(16'hffff);
  assign T6447 = {T6450, T6448};
  assign T6448 = $signed(T6449) / $signed(22'h100000);
  assign T6449 = $signed(30'h24a2eff7) * $signed(16'h0);
  assign T6450 = T6448[6'h2d:6'h2d];
  assign twiddle4_3_465_imag = T6453 + T6451;
  assign T6451 = $signed(T6452) / $signed(22'h100000);
  assign T6452 = $signed(31'h45e531a2) * $signed(16'hffff);
  assign T6453 = {T6456, T6454};
  assign T6454 = $signed(T6455) / $signed(22'h100000);
  assign T6455 = $signed(30'h252b8cee) * $signed(16'h0);
  assign T6456 = T6454[6'h2d:6'h2d];
  assign T6457 = T2943[1'h0:1'h0];
  assign T6458 = T6471 ? twiddle4_3_467_imag : twiddle4_3_466_imag;
  assign twiddle4_3_466_imag = T6461 + T6459;
  assign T6459 = $signed(T6460) / $signed(22'h100000);
  assign T6460 = $signed(31'h45a69bbf) * $signed(16'hffff);
  assign T6461 = {T6464, T6462};
  assign T6462 = $signed(T6463) / $signed(22'h100000);
  assign T6463 = $signed(30'h25b4bed9) * $signed(16'h0);
  assign T6464 = T6462[6'h2d:6'h2d];
  assign twiddle4_3_467_imag = T6467 + T6465;
  assign T6465 = $signed(T6466) / $signed(22'h100000);
  assign T6466 = $signed(31'h456949ca) * $signed(16'hffff);
  assign T6467 = {T6470, T6468};
  assign T6468 = $signed(T6469) / $signed(22'h100000);
  assign T6469 = $signed(30'h263e82bc) * $signed(16'h0);
  assign T6470 = T6468[6'h2d:6'h2d];
  assign T6471 = T2943[1'h0:1'h0];
  assign T6472 = T2943[1'h1:1'h1];
  assign T6473 = T6502 ? T6488 : T6474;
  assign T6474 = T6487 ? twiddle4_3_469_imag : twiddle4_3_468_imag;
  assign twiddle4_3_468_imag = T6477 + T6475;
  assign T6475 = $signed(T6476) / $signed(22'h100000);
  assign T6476 = $signed(31'h452d3d19) * $signed(16'hffff);
  assign T6477 = {T6480, T6478};
  assign T6478 = $signed(T6479) / $signed(22'h100000);
  assign T6479 = $signed(30'h26c8d59d) * $signed(16'h0);
  assign T6480 = T6478[6'h2d:6'h2d];
  assign twiddle4_3_469_imag = T6483 + T6481;
  assign T6481 = $signed(T6482) / $signed(22'h100000);
  assign T6482 = $signed(31'h44f276f8) * $signed(16'hffff);
  assign T6483 = {T6486, T6484};
  assign T6484 = $signed(T6485) / $signed(22'h100000);
  assign T6485 = $signed(30'h2753b47a) * $signed(16'h0);
  assign T6486 = T6484[6'h2d:6'h2d];
  assign T6487 = T2943[1'h0:1'h0];
  assign T6488 = T6501 ? twiddle4_3_471_imag : twiddle4_3_470_imag;
  assign twiddle4_3_470_imag = T6491 + T6489;
  assign T6489 = $signed(T6490) / $signed(22'h100000);
  assign T6490 = $signed(31'h44b8f8ae) * $signed(16'hffff);
  assign T6491 = {T6494, T6492};
  assign T6492 = $signed(T6493) / $signed(22'h100000);
  assign T6493 = $signed(30'h27df1c50) * $signed(16'h0);
  assign T6494 = T6492[6'h2d:6'h2d];
  assign twiddle4_3_471_imag = T6497 + T6495;
  assign T6495 = $signed(T6496) / $signed(22'h100000);
  assign T6496 = $signed(31'h4480c379) * $signed(16'hffff);
  assign T6497 = {T6500, T6498};
  assign T6498 = $signed(T6499) / $signed(22'h100000);
  assign T6499 = $signed(30'h286b0a1a) * $signed(16'h0);
  assign T6500 = T6498[6'h2d:6'h2d];
  assign T6501 = T2943[1'h0:1'h0];
  assign T6502 = T2943[1'h1:1'h1];
  assign T6503 = T2943[2'h2:2'h2];
  assign T6504 = T6565 ? T6535 : T6505;
  assign T6505 = T6534 ? T6520 : T6506;
  assign T6506 = T6519 ? twiddle4_3_473_imag : twiddle4_3_472_imag;
  assign twiddle4_3_472_imag = T6509 + T6507;
  assign T6507 = $signed(T6508) / $signed(22'h100000);
  assign T6508 = $signed(31'h4449d893) * $signed(16'hffff);
  assign T6509 = {T6512, T6510};
  assign T6510 = $signed(T6511) / $signed(22'h100000);
  assign T6511 = $signed(30'h28f77ad0) * $signed(16'h0);
  assign T6512 = T6510[6'h2d:6'h2d];
  assign twiddle4_3_473_imag = T6515 + T6513;
  assign T6513 = $signed(T6514) / $signed(22'h100000);
  assign T6514 = $signed(31'h4414392b) * $signed(16'hffff);
  assign T6515 = {T6518, T6516};
  assign T6516 = $signed(T6517) / $signed(22'h100000);
  assign T6517 = $signed(30'h29846b64) * $signed(16'h0);
  assign T6518 = T6516[6'h2d:6'h2d];
  assign T6519 = T2943[1'h0:1'h0];
  assign T6520 = T6533 ? twiddle4_3_475_imag : twiddle4_3_474_imag;
  assign twiddle4_3_474_imag = T6523 + T6521;
  assign T6521 = $signed(T6522) / $signed(22'h100000);
  assign T6522 = $signed(31'h43dfe66c) * $signed(16'hffff);
  assign T6523 = {T6526, T6524};
  assign T6524 = $signed(T6525) / $signed(22'h100000);
  assign T6525 = $signed(30'h2a11d8c9) * $signed(16'h0);
  assign T6526 = T6524[6'h2d:6'h2d];
  assign twiddle4_3_475_imag = T6529 + T6527;
  assign T6527 = $signed(T6528) / $signed(22'h100000);
  assign T6528 = $signed(31'h43ace178) * $signed(16'hffff);
  assign T6529 = {T6532, T6530};
  assign T6530 = $signed(T6531) / $signed(22'h100000);
  assign T6531 = $signed(30'h2a9fbfee) * $signed(16'h0);
  assign T6532 = T6530[6'h2d:6'h2d];
  assign T6533 = T2943[1'h0:1'h0];
  assign T6534 = T2943[1'h1:1'h1];
  assign T6535 = T6564 ? T6550 : T6536;
  assign T6536 = T6549 ? twiddle4_3_477_imag : twiddle4_3_476_imag;
  assign twiddle4_3_476_imag = T6539 + T6537;
  assign T6537 = $signed(T6538) / $signed(22'h100000);
  assign T6538 = $signed(31'h437b2b6a) * $signed(16'hffff);
  assign T6539 = {T6542, T6540};
  assign T6540 = $signed(T6541) / $signed(22'h100000);
  assign T6541 = $signed(30'h2b2e1dbe) * $signed(16'h0);
  assign T6542 = T6540[6'h2d:6'h2d];
  assign twiddle4_3_477_imag = T6545 + T6543;
  assign T6543 = $signed(T6544) / $signed(22'h100000);
  assign T6544 = $signed(31'h434ac556) * $signed(16'hffff);
  assign T6545 = {T6548, T6546};
  assign T6546 = $signed(T6547) / $signed(22'h100000);
  assign T6547 = $signed(30'h2bbcef24) * $signed(16'h0);
  assign T6548 = T6546[6'h2d:6'h2d];
  assign T6549 = T2943[1'h0:1'h0];
  assign T6550 = T6563 ? twiddle4_3_479_imag : twiddle4_3_478_imag;
  assign twiddle4_3_478_imag = T6553 + T6551;
  assign T6551 = $signed(T6552) / $signed(22'h100000);
  assign T6552 = $signed(31'h431bb04a) * $signed(16'hffff);
  assign T6553 = {T6556, T6554};
  assign T6554 = $signed(T6555) / $signed(22'h100000);
  assign T6555 = $signed(30'h2c4c3106) * $signed(16'h0);
  assign T6556 = T6554[6'h2d:6'h2d];
  assign twiddle4_3_479_imag = T6559 + T6557;
  assign T6557 = $signed(T6558) / $signed(22'h100000);
  assign T6558 = $signed(31'h42eded49) * $signed(16'hffff);
  assign T6559 = {T6562, T6560};
  assign T6560 = $signed(T6561) / $signed(22'h100000);
  assign T6561 = $signed(30'h2cdbe04a) * $signed(16'h0);
  assign T6562 = T6560[6'h2d:6'h2d];
  assign T6563 = T2943[1'h0:1'h0];
  assign T6564 = T2943[1'h1:1'h1];
  assign T6565 = T2943[2'h2:2'h2];
  assign T6566 = T2943[2'h3:2'h3];
  assign T6567 = T2943[3'h4:3'h4];
  assign T6568 = T6848 ? T6706 : T6569;
  assign T6569 = T6705 ? T6635 : T6570;
  assign T6570 = T6634 ? T6601 : T6571;
  assign T6571 = T6600 ? T6586 : T6572;
  assign T6572 = T6585 ? twiddle4_3_481_imag : twiddle4_3_480_imag;
  assign twiddle4_3_480_imag = T6575 + T6573;
  assign T6573 = $signed(T6574) / $signed(22'h100000);
  assign T6574 = $signed(31'h42c17d53) * $signed(16'hffff);
  assign T6575 = {T6578, T6576};
  assign T6576 = $signed(T6577) / $signed(22'h100000);
  assign T6577 = $signed(30'h2d6bf9d2) * $signed(16'h0);
  assign T6578 = T6576[6'h2d:6'h2d];
  assign twiddle4_3_481_imag = T6581 + T6579;
  assign T6579 = $signed(T6580) / $signed(22'h100000);
  assign T6580 = $signed(31'h4296615e) * $signed(16'hffff);
  assign T6581 = {T6584, T6582};
  assign T6582 = $signed(T6583) / $signed(22'h100000);
  assign T6583 = $signed(30'h2dfc7a7d) * $signed(16'h0);
  assign T6584 = T6582[6'h2d:6'h2d];
  assign T6585 = T2943[1'h0:1'h0];
  assign T6586 = T6599 ? twiddle4_3_483_imag : twiddle4_3_482_imag;
  assign twiddle4_3_482_imag = T6589 + T6587;
  assign T6587 = $signed(T6588) / $signed(22'h100000);
  assign T6588 = $signed(31'h426c9a59) * $signed(16'hffff);
  assign T6589 = {T6592, T6590};
  assign T6590 = $signed(T6591) / $signed(22'h100000);
  assign T6591 = $signed(30'h2e8d5f29) * $signed(16'h0);
  assign T6592 = T6590[6'h2d:6'h2d];
  assign twiddle4_3_483_imag = T6595 + T6593;
  assign T6593 = $signed(T6594) / $signed(22'h100000);
  assign T6594 = $signed(31'h4244292c) * $signed(16'hffff);
  assign T6595 = {T6598, T6596};
  assign T6596 = $signed(T6597) / $signed(22'h100000);
  assign T6597 = $signed(30'h2f1ea4b2) * $signed(16'h0);
  assign T6598 = T6596[6'h2d:6'h2d];
  assign T6599 = T2943[1'h0:1'h0];
  assign T6600 = T2943[1'h1:1'h1];
  assign T6601 = T6633 ? T6617 : T6602;
  assign T6602 = T6616 ? twiddle4_3_485_imag : twiddle4_3_484_imag;
  assign twiddle4_3_484_imag = T6605 + T6603;
  assign T6603 = $signed(T6604) / $signed(22'h100000);
  assign T6604 = $signed(31'h421d0eb9) * $signed(16'hffff);
  assign T6605 = {T6608, T6606};
  assign T6606 = $signed(T6607) / $signed(22'h100000);
  assign T6607 = $signed(30'h2fb047f2) * $signed(16'h0);
  assign T6608 = T6606[6'h2d:6'h2d];
  assign twiddle4_3_485_imag = T6611 + T6609;
  assign T6609 = $signed(T6610) / $signed(22'h100000);
  assign T6610 = $signed(31'h41f74bd7) * $signed(16'hffff);
  assign T6611 = {T6614, T6612};
  assign T6612 = $signed(T6613) / $signed(22'h100000);
  assign T6613 = $signed(29'h104245c0) * $signed(16'h0);
  assign T6614 = T6615 ? 2'h3 : 2'h0;
  assign T6615 = T6612[6'h2c:6'h2c];
  assign T6616 = T2943[1'h0:1'h0];
  assign T6617 = T6632 ? twiddle4_3_487_imag : twiddle4_3_486_imag;
  assign twiddle4_3_486_imag = T6620 + T6618;
  assign T6618 = $signed(T6619) / $signed(22'h100000);
  assign T6619 = $signed(31'h41d2e159) * $signed(16'hffff);
  assign T6620 = {T6623, T6621};
  assign T6621 = $signed(T6622) / $signed(22'h100000);
  assign T6622 = $signed(29'h10d49af1) * $signed(16'h0);
  assign T6623 = T6624 ? 2'h3 : 2'h0;
  assign T6624 = T6621[6'h2c:6'h2c];
  assign twiddle4_3_487_imag = T6627 + T6625;
  assign T6625 = $signed(T6626) / $signed(22'h100000);
  assign T6626 = $signed(31'h41afd008) * $signed(16'hffff);
  assign T6627 = {T6630, T6628};
  assign T6628 = $signed(T6629) / $signed(22'h100000);
  assign T6629 = $signed(29'h1167445a) * $signed(16'h0);
  assign T6630 = T6631 ? 2'h3 : 2'h0;
  assign T6631 = T6628[6'h2c:6'h2c];
  assign T6632 = T2943[1'h0:1'h0];
  assign T6633 = T2943[1'h1:1'h1];
  assign T6634 = T2943[2'h2:2'h2];
  assign T6635 = T6704 ? T6670 : T6636;
  assign T6636 = T6669 ? T6653 : T6637;
  assign T6637 = T6652 ? twiddle4_3_489_imag : twiddle4_3_488_imag;
  assign twiddle4_3_488_imag = T6640 + T6638;
  assign T6638 = $signed(T6639) / $signed(22'h100000);
  assign T6639 = $signed(31'h418e18a8) * $signed(16'hffff);
  assign T6640 = {T6643, T6641};
  assign T6641 = $signed(T6642) / $signed(22'h100000);
  assign T6642 = $signed(29'h11fa3ecb) * $signed(16'h0);
  assign T6643 = T6644 ? 2'h3 : 2'h0;
  assign T6644 = T6641[6'h2c:6'h2c];
  assign twiddle4_3_489_imag = T6647 + T6645;
  assign T6645 = $signed(T6646) / $signed(22'h100000);
  assign T6646 = $signed(31'h416dbbf3) * $signed(16'hffff);
  assign T6647 = {T6650, T6648};
  assign T6648 = $signed(T6649) / $signed(22'h100000);
  assign T6649 = $signed(29'h128d8716) * $signed(16'h0);
  assign T6650 = T6651 ? 2'h3 : 2'h0;
  assign T6651 = T6648[6'h2c:6'h2c];
  assign T6652 = T2943[1'h0:1'h0];
  assign T6653 = T6668 ? twiddle4_3_491_imag : twiddle4_3_490_imag;
  assign twiddle4_3_490_imag = T6656 + T6654;
  assign T6654 = $signed(T6655) / $signed(22'h100000);
  assign T6655 = $signed(31'h414eba9e) * $signed(16'hffff);
  assign T6656 = {T6659, T6657};
  assign T6657 = $signed(T6658) / $signed(22'h100000);
  assign T6658 = $signed(29'h13211a07) * $signed(16'h0);
  assign T6659 = T6660 ? 2'h3 : 2'h0;
  assign T6660 = T6657[6'h2c:6'h2c];
  assign twiddle4_3_491_imag = T6663 + T6661;
  assign T6661 = $signed(T6662) / $signed(22'h100000);
  assign T6662 = $signed(31'h41311553) * $signed(16'hffff);
  assign T6663 = {T6666, T6664};
  assign T6664 = $signed(T6665) / $signed(22'h100000);
  assign T6665 = $signed(29'h13b4f46d) * $signed(16'h0);
  assign T6666 = T6667 ? 2'h3 : 2'h0;
  assign T6667 = T6664[6'h2c:6'h2c];
  assign T6668 = T2943[1'h0:1'h0];
  assign T6669 = T2943[1'h1:1'h1];
  assign T6670 = T6703 ? T6687 : T6671;
  assign T6671 = T6686 ? twiddle4_3_493_imag : twiddle4_3_492_imag;
  assign twiddle4_3_492_imag = T6674 + T6672;
  assign T6672 = $signed(T6673) / $signed(22'h100000);
  assign T6673 = $signed(31'h4114ccb9) * $signed(16'hffff);
  assign T6674 = {T6677, T6675};
  assign T6675 = $signed(T6676) / $signed(22'h100000);
  assign T6676 = $signed(29'h14491311) * $signed(16'h0);
  assign T6677 = T6678 ? 2'h3 : 2'h0;
  assign T6678 = T6675[6'h2c:6'h2c];
  assign twiddle4_3_493_imag = T6681 + T6679;
  assign T6679 = $signed(T6680) / $signed(22'h100000);
  assign T6680 = $signed(31'h40f9e16c) * $signed(16'hffff);
  assign T6681 = {T6684, T6682};
  assign T6682 = $signed(T6683) / $signed(22'h100000);
  assign T6683 = $signed(29'h14dd72bf) * $signed(16'h0);
  assign T6684 = T6685 ? 2'h3 : 2'h0;
  assign T6685 = T6682[6'h2c:6'h2c];
  assign T6686 = T2943[1'h0:1'h0];
  assign T6687 = T6702 ? twiddle4_3_495_imag : twiddle4_3_494_imag;
  assign twiddle4_3_494_imag = T6690 + T6688;
  assign T6688 = $signed(T6689) / $signed(22'h100000);
  assign T6689 = $signed(31'h40e05401) * $signed(16'hffff);
  assign T6690 = {T6693, T6691};
  assign T6691 = $signed(T6692) / $signed(22'h100000);
  assign T6692 = $signed(29'h1572103e) * $signed(16'h0);
  assign T6693 = T6694 ? 2'h3 : 2'h0;
  assign T6694 = T6691[6'h2c:6'h2c];
  assign twiddle4_3_495_imag = T6697 + T6695;
  assign T6695 = $signed(T6696) / $signed(22'h100000);
  assign T6696 = $signed(31'h40c82507) * $signed(16'hffff);
  assign T6697 = {T6700, T6698};
  assign T6698 = $signed(T6699) / $signed(22'h100000);
  assign T6699 = $signed(29'h1606e855) * $signed(16'h0);
  assign T6700 = T6701 ? 2'h3 : 2'h0;
  assign T6701 = T6698[6'h2c:6'h2c];
  assign T6702 = T2943[1'h0:1'h0];
  assign T6703 = T2943[1'h1:1'h1];
  assign T6704 = T2943[2'h2:2'h2];
  assign T6705 = T2943[2'h3:2'h3];
  assign T6706 = T6847 ? T6777 : T6707;
  assign T6707 = T6776 ? T6742 : T6708;
  assign T6708 = T6741 ? T6725 : T6709;
  assign T6709 = T6724 ? twiddle4_3_497_imag : twiddle4_3_496_imag;
  assign twiddle4_3_496_imag = T6712 + T6710;
  assign T6710 = $signed(T6711) / $signed(22'h100000);
  assign T6711 = $signed(31'h40b15502) * $signed(16'hffff);
  assign T6712 = {T6715, T6713};
  assign T6713 = $signed(T6714) / $signed(22'h100000);
  assign T6714 = $signed(29'h169bf7c9) * $signed(16'h0);
  assign T6715 = T6716 ? 2'h3 : 2'h0;
  assign T6716 = T6713[6'h2c:6'h2c];
  assign twiddle4_3_497_imag = T6719 + T6717;
  assign T6717 = $signed(T6718) / $signed(22'h100000);
  assign T6718 = $signed(31'h409be473) * $signed(16'hffff);
  assign T6719 = {T6722, T6720};
  assign T6720 = $signed(T6721) / $signed(22'h100000);
  assign T6721 = $signed(29'h17313b60) * $signed(16'h0);
  assign T6722 = T6723 ? 2'h3 : 2'h0;
  assign T6723 = T6720[6'h2c:6'h2c];
  assign T6724 = T2943[1'h0:1'h0];
  assign T6725 = T6740 ? twiddle4_3_499_imag : twiddle4_3_498_imag;
  assign twiddle4_3_498_imag = T6728 + T6726;
  assign T6726 = $signed(T6727) / $signed(22'h100000);
  assign T6727 = $signed(31'h4087d3d1) * $signed(16'hffff);
  assign T6728 = {T6731, T6729};
  assign T6729 = $signed(T6730) / $signed(22'h100000);
  assign T6730 = $signed(29'h17c6afdd) * $signed(16'h0);
  assign T6731 = T6732 ? 2'h3 : 2'h0;
  assign T6732 = T6729[6'h2c:6'h2c];
  assign twiddle4_3_499_imag = T6735 + T6733;
  assign T6733 = $signed(T6734) / $signed(22'h100000);
  assign T6734 = $signed(31'h4075238a) * $signed(16'hffff);
  assign T6735 = {T6738, T6736};
  assign T6736 = $signed(T6737) / $signed(22'h100000);
  assign T6737 = $signed(28'h85c5201) * $signed(16'h0);
  assign T6738 = T6739 ? 3'h7 : 3'h0;
  assign T6739 = T6736[6'h2b:6'h2b];
  assign T6740 = T2943[1'h0:1'h0];
  assign T6741 = T2943[1'h1:1'h1];
  assign T6742 = T6775 ? T6759 : T6743;
  assign T6743 = T6758 ? twiddle4_3_501_imag : twiddle4_3_500_imag;
  assign twiddle4_3_500_imag = T6746 + T6744;
  assign T6744 = $signed(T6745) / $signed(22'h100000);
  assign T6745 = $signed(31'h4063d406) * $signed(16'hffff);
  assign T6746 = {T6749, T6747};
  assign T6747 = $signed(T6748) / $signed(22'h100000);
  assign T6748 = $signed(28'h8f21e8f) * $signed(16'h0);
  assign T6749 = T6750 ? 3'h7 : 3'h0;
  assign T6750 = T6747[6'h2b:6'h2b];
  assign twiddle4_3_501_imag = T6753 + T6751;
  assign T6751 = $signed(T6752) / $signed(22'h100000);
  assign T6752 = $signed(31'h4053e5a5) * $signed(16'hffff);
  assign T6753 = {T6756, T6754};
  assign T6754 = $signed(T6755) / $signed(22'h100000);
  assign T6755 = $signed(28'h9881246) * $signed(16'h0);
  assign T6756 = T6757 ? 3'h7 : 3'h0;
  assign T6757 = T6754[6'h2b:6'h2b];
  assign T6758 = T2943[1'h0:1'h0];
  assign T6759 = T6774 ? twiddle4_3_503_imag : twiddle4_3_502_imag;
  assign twiddle4_3_502_imag = T6762 + T6760;
  assign T6760 = $signed(T6761) / $signed(22'h100000);
  assign T6761 = $signed(31'h404558c1) * $signed(16'hffff);
  assign T6762 = {T6765, T6763};
  assign T6763 = $signed(T6764) / $signed(22'h100000);
  assign T6764 = $signed(28'ha1e29e6) * $signed(16'h0);
  assign T6765 = T6766 ? 3'h7 : 3'h0;
  assign T6766 = T6763[6'h2b:6'h2b];
  assign twiddle4_3_503_imag = T6769 + T6767;
  assign T6767 = $signed(T6768) / $signed(22'h100000);
  assign T6768 = $signed(31'h40382da9) * $signed(16'hffff);
  assign T6769 = {T6772, T6770};
  assign T6770 = $signed(T6771) / $signed(22'h100000);
  assign T6771 = $signed(28'hab4622e) * $signed(16'h0);
  assign T6772 = T6773 ? 3'h7 : 3'h0;
  assign T6773 = T6770[6'h2b:6'h2b];
  assign T6774 = T2943[1'h0:1'h0];
  assign T6775 = T2943[1'h1:1'h1];
  assign T6776 = T2943[2'h2:2'h2];
  assign T6777 = T6846 ? T6812 : T6778;
  assign T6778 = T6811 ? T6795 : T6779;
  assign T6779 = T6794 ? twiddle4_3_505_imag : twiddle4_3_504_imag;
  assign twiddle4_3_504_imag = T6782 + T6780;
  assign T6780 = $signed(T6781) / $signed(22'h100000);
  assign T6781 = $signed(31'h402c64a6) * $signed(16'hffff);
  assign T6782 = {T6785, T6783};
  assign T6783 = $signed(T6784) / $signed(22'h100000);
  assign T6784 = $signed(28'hb4ab7dc) * $signed(16'h0);
  assign T6785 = T6786 ? 3'h7 : 3'h0;
  assign T6786 = T6783[6'h2b:6'h2b];
  assign twiddle4_3_505_imag = T6789 + T6787;
  assign T6787 = $signed(T6788) / $signed(22'h100000);
  assign T6788 = $signed(31'h4021fdfb) * $signed(16'hffff);
  assign T6789 = {T6792, T6790};
  assign T6790 = $signed(T6791) / $signed(22'h100000);
  assign T6791 = $signed(28'hbe127ad) * $signed(16'h0);
  assign T6792 = T6793 ? 3'h7 : 3'h0;
  assign T6793 = T6790[6'h2b:6'h2b];
  assign T6794 = T2943[1'h0:1'h0];
  assign T6795 = T6810 ? twiddle4_3_507_imag : twiddle4_3_506_imag;
  assign twiddle4_3_506_imag = T6798 + T6796;
  assign T6796 = $signed(T6797) / $signed(22'h100000);
  assign T6797 = $signed(31'h4018f9e1) * $signed(16'hffff);
  assign T6798 = {T6801, T6799};
  assign T6799 = $signed(T6800) / $signed(22'h100000);
  assign T6800 = $signed(27'h477ae5e) * $signed(16'h0);
  assign T6801 = T6802 ? 4'hf : 4'h0;
  assign T6802 = T6799[6'h2a:6'h2a];
  assign twiddle4_3_507_imag = T6805 + T6803;
  assign T6803 = $signed(T6804) / $signed(22'h100000);
  assign T6804 = $signed(31'h4011588a) * $signed(16'hffff);
  assign T6805 = {T6808, T6806};
  assign T6806 = $signed(T6807) / $signed(22'h100000);
  assign T6807 = $signed(27'h50e48ac) * $signed(16'h0);
  assign T6808 = T6809 ? 4'hf : 4'h0;
  assign T6809 = T6806[6'h2a:6'h2a];
  assign T6810 = T2943[1'h0:1'h0];
  assign T6811 = T2943[1'h1:1'h1];
  assign T6812 = T6845 ? T6829 : T6813;
  assign T6813 = T6828 ? twiddle4_3_509_imag : twiddle4_3_508_imag;
  assign twiddle4_3_508_imag = T6816 + T6814;
  assign T6814 = $signed(T6815) / $signed(22'h100000);
  assign T6815 = $signed(31'h400b1a21) * $signed(16'hffff);
  assign T6816 = {T6819, T6817};
  assign T6817 = $signed(T6818) / $signed(22'h100000);
  assign T6818 = $signed(27'h5a4f352) * $signed(16'h0);
  assign T6819 = T6820 ? 4'hf : 4'h0;
  assign T6820 = T6817[6'h2a:6'h2a];
  assign twiddle4_3_509_imag = T6823 + T6821;
  assign T6821 = $signed(T6822) / $signed(22'h100000);
  assign T6822 = $signed(31'h40063ec7) * $signed(16'hffff);
  assign T6823 = {T6826, T6824};
  assign T6824 = $signed(T6825) / $signed(22'h100000);
  assign T6825 = $signed(26'h23bab0c) * $signed(16'h0);
  assign T6826 = T6827 ? 5'h1f : 5'h0;
  assign T6827 = T6824[6'h29:6'h29];
  assign T6828 = T2943[1'h0:1'h0];
  assign T6829 = T6844 ? twiddle4_3_511_imag : twiddle4_3_510_imag;
  assign twiddle4_3_510_imag = T6832 + T6830;
  assign T6830 = $signed(T6831) / $signed(22'h100000);
  assign T6831 = $signed(31'h4002c698) * $signed(16'hffff);
  assign T6832 = {T6835, T6833};
  assign T6833 = $signed(T6834) / $signed(22'h100000);
  assign T6834 = $signed(26'h2d26c95) * $signed(16'h0);
  assign T6835 = T6836 ? 5'h1f : 5'h0;
  assign T6836 = T6833[6'h29:6'h29];
  assign twiddle4_3_511_imag = T6839 + T6837;
  assign T6837 = $signed(T6838) / $signed(22'h100000);
  assign T6838 = $signed(31'h4000b1a7) * $signed(16'hffff);
  assign T6839 = {T6842, T6840};
  assign T6840 = $signed(T6841) / $signed(22'h100000);
  assign T6841 = $signed(25'h16934a8) * $signed(16'h0);
  assign T6842 = T6843 ? 6'h3f : 6'h0;
  assign T6843 = T6840[6'h28:6'h28];
  assign T6844 = T2943[1'h0:1'h0];
  assign T6845 = T2943[1'h1:1'h1];
  assign T6846 = T2943[2'h2:2'h2];
  assign T6847 = T2943[2'h3:2'h3];
  assign T6848 = T2943[3'h4:3'h4];
  assign T6849 = T2943[3'h5:3'h5];
  assign T6850 = T2943[3'h6:3'h6];
  assign T6851 = T2943[3'h7:3'h7];
  assign T6852 = T4896[6'h2e:6'h2e];
  assign T6853 = T2943[4'h8:4'h8];
  assign io_t4_3out_real = T6854;
  assign T6854 = T6855[4'hf:1'h0];
  assign T6855 = T10789 ? T8831 : T6856;
  assign T6856 = T8830 ? T7807 : T6857;
  assign T6857 = T7806 ? T7394 : T6858;
  assign T6858 = T7393 ? T7151 : T6859;
  assign T6859 = T7150 ? T7010 : T6860;
  assign T6860 = T7009 ? T6937 : T6861;
  assign T6861 = T6936 ? T6900 : T6862;
  assign T6862 = T6899 ? T6881 : T6863;
  assign T6863 = T6880 ? T6871 : twiddle4_3_0_real;
  assign twiddle4_3_0_real = T6869 + T6864;
  assign T6864 = {T6867, T6865};
  assign T6865 = $signed(T6866) / $signed(22'h100000);
  assign T6866 = $signed(1'h0) * $signed(16'h0);
  assign T6867 = T6868 ? 31'h7fffffff : 31'h0;
  assign T6868 = T6865[5'h10:5'h10];
  assign T6869 = $signed(T6870) / $signed(22'h100000);
  assign T6870 = $signed(32'h40000000) * $signed(16'h1);
  assign T6871 = {T6879, twiddle4_3_1_real};
  assign twiddle4_3_1_real = T6877 + T6872;
  assign T6872 = {T6875, T6873};
  assign T6873 = $signed(T6874) / $signed(22'h100000);
  assign T6874 = $signed(25'h96cb58) * $signed(16'h0);
  assign T6875 = T6876 ? 6'h3f : 6'h0;
  assign T6876 = T6873[6'h28:6'h28];
  assign T6877 = $signed(T6878) / $signed(22'h100000);
  assign T6878 = $signed(31'h3fff4e59) * $signed(16'h1);
  assign T6879 = twiddle4_3_1_real[6'h2e:6'h2e];
  assign T6880 = T2943[1'h0:1'h0];
  assign T6881 = {T6898, T6882};
  assign T6882 = T6897 ? twiddle4_3_3_real : twiddle4_3_2_real;
  assign twiddle4_3_2_real = T6888 + T6883;
  assign T6883 = {T6886, T6884};
  assign T6884 = $signed(T6885) / $signed(22'h100000);
  assign T6885 = $signed(26'h12d936b) * $signed(16'h0);
  assign T6886 = T6887 ? 5'h1f : 5'h0;
  assign T6887 = T6884[6'h29:6'h29];
  assign T6888 = $signed(T6889) / $signed(22'h100000);
  assign T6889 = $signed(31'h3ffd3968) * $signed(16'h1);
  assign twiddle4_3_3_real = T6895 + T6890;
  assign T6890 = {T6893, T6891};
  assign T6891 = $signed(T6892) / $signed(22'h100000);
  assign T6892 = $signed(26'h1c454f4) * $signed(16'h0);
  assign T6893 = T6894 ? 5'h1f : 5'h0;
  assign T6894 = T6891[6'h29:6'h29];
  assign T6895 = $signed(T6896) / $signed(22'h100000);
  assign T6896 = $signed(31'h3ff9c139) * $signed(16'h1);
  assign T6897 = T2943[1'h0:1'h0];
  assign T6898 = T6882[6'h2e:6'h2e];
  assign T6899 = T2943[1'h1:1'h1];
  assign T6900 = {T6935, T6901};
  assign T6901 = T6934 ? T6918 : T6902;
  assign T6902 = T6917 ? twiddle4_3_5_real : twiddle4_3_4_real;
  assign twiddle4_3_4_real = T6908 + T6903;
  assign T6903 = {T6906, T6904};
  assign T6904 = $signed(T6905) / $signed(22'h100000);
  assign T6905 = $signed(27'h25b0cae) * $signed(16'h0);
  assign T6906 = T6907 ? 4'hf : 4'h0;
  assign T6907 = T6904[6'h2a:6'h2a];
  assign T6908 = $signed(T6909) / $signed(22'h100000);
  assign T6909 = $signed(31'h3ff4e5df) * $signed(16'h1);
  assign twiddle4_3_5_real = T6915 + T6910;
  assign T6910 = {T6913, T6911};
  assign T6911 = $signed(T6912) / $signed(22'h100000);
  assign T6912 = $signed(27'h2f1b754) * $signed(16'h0);
  assign T6913 = T6914 ? 4'hf : 4'h0;
  assign T6914 = T6911[6'h2a:6'h2a];
  assign T6915 = $signed(T6916) / $signed(22'h100000);
  assign T6916 = $signed(31'h3feea776) * $signed(16'h1);
  assign T6917 = T2943[1'h0:1'h0];
  assign T6918 = T6933 ? twiddle4_3_7_real : twiddle4_3_6_real;
  assign twiddle4_3_6_real = T6924 + T6919;
  assign T6919 = {T6922, T6920};
  assign T6920 = $signed(T6921) / $signed(22'h100000);
  assign T6921 = $signed(27'h38851a2) * $signed(16'h0);
  assign T6922 = T6923 ? 4'hf : 4'h0;
  assign T6923 = T6920[6'h2a:6'h2a];
  assign T6924 = $signed(T6925) / $signed(22'h100000);
  assign T6925 = $signed(31'h3fe7061f) * $signed(16'h1);
  assign twiddle4_3_7_real = T6931 + T6926;
  assign T6926 = {T6929, T6927};
  assign T6927 = $signed(T6928) / $signed(22'h100000);
  assign T6928 = $signed(28'h41ed853) * $signed(16'h0);
  assign T6929 = T6930 ? 3'h7 : 3'h0;
  assign T6930 = T6927[6'h2b:6'h2b];
  assign T6931 = $signed(T6932) / $signed(22'h100000);
  assign T6932 = $signed(31'h3fde0205) * $signed(16'h1);
  assign T6933 = T2943[1'h0:1'h0];
  assign T6934 = T2943[1'h1:1'h1];
  assign T6935 = T6901[6'h2e:6'h2e];
  assign T6936 = T2943[2'h2:2'h2];
  assign T6937 = {T7008, T6938};
  assign T6938 = T7007 ? T6973 : T6939;
  assign T6939 = T6972 ? T6956 : T6940;
  assign T6940 = T6955 ? twiddle4_3_9_real : twiddle4_3_8_real;
  assign twiddle4_3_8_real = T6946 + T6941;
  assign T6941 = {T6944, T6942};
  assign T6942 = $signed(T6943) / $signed(22'h100000);
  assign T6943 = $signed(28'h4b54824) * $signed(16'h0);
  assign T6944 = T6945 ? 3'h7 : 3'h0;
  assign T6945 = T6942[6'h2b:6'h2b];
  assign T6946 = $signed(T6947) / $signed(22'h100000);
  assign T6947 = $signed(31'h3fd39b5a) * $signed(16'h1);
  assign twiddle4_3_9_real = T6953 + T6948;
  assign T6948 = {T6951, T6949};
  assign T6949 = $signed(T6950) / $signed(22'h100000);
  assign T6950 = $signed(28'h54b9dd2) * $signed(16'h0);
  assign T6951 = T6952 ? 3'h7 : 3'h0;
  assign T6952 = T6949[6'h2b:6'h2b];
  assign T6953 = $signed(T6954) / $signed(22'h100000);
  assign T6954 = $signed(31'h3fc7d257) * $signed(16'h1);
  assign T6955 = T2943[1'h0:1'h0];
  assign T6956 = T6971 ? twiddle4_3_11_real : twiddle4_3_10_real;
  assign twiddle4_3_10_real = T6962 + T6957;
  assign T6957 = {T6960, T6958};
  assign T6958 = $signed(T6959) / $signed(22'h100000);
  assign T6959 = $signed(28'h5e1d61a) * $signed(16'h0);
  assign T6960 = T6961 ? 3'h7 : 3'h0;
  assign T6961 = T6958[6'h2b:6'h2b];
  assign T6962 = $signed(T6963) / $signed(22'h100000);
  assign T6963 = $signed(31'h3fbaa73f) * $signed(16'h1);
  assign twiddle4_3_11_real = T6969 + T6964;
  assign T6964 = {T6967, T6965};
  assign T6965 = $signed(T6966) / $signed(22'h100000);
  assign T6966 = $signed(28'h677edba) * $signed(16'h0);
  assign T6967 = T6968 ? 3'h7 : 3'h0;
  assign T6968 = T6965[6'h2b:6'h2b];
  assign T6969 = $signed(T6970) / $signed(22'h100000);
  assign T6970 = $signed(31'h3fac1a5b) * $signed(16'h1);
  assign T6971 = T2943[1'h0:1'h0];
  assign T6972 = T2943[1'h1:1'h1];
  assign T6973 = T7006 ? T6990 : T6974;
  assign T6974 = T6989 ? twiddle4_3_13_real : twiddle4_3_12_real;
  assign twiddle4_3_12_real = T6980 + T6975;
  assign T6975 = {T6978, T6976};
  assign T6976 = $signed(T6977) / $signed(22'h100000);
  assign T6977 = $signed(28'h70de171) * $signed(16'h0);
  assign T6978 = T6979 ? 3'h7 : 3'h0;
  assign T6979 = T6976[6'h2b:6'h2b];
  assign T6980 = $signed(T6981) / $signed(22'h100000);
  assign T6981 = $signed(31'h3f9c2bfa) * $signed(16'h1);
  assign twiddle4_3_13_real = T6987 + T6982;
  assign T6982 = {T6985, T6983};
  assign T6983 = $signed(T6984) / $signed(22'h100000);
  assign T6984 = $signed(28'h7a3adff) * $signed(16'h0);
  assign T6985 = T6986 ? 3'h7 : 3'h0;
  assign T6986 = T6983[6'h2b:6'h2b];
  assign T6987 = $signed(T6988) / $signed(22'h100000);
  assign T6988 = $signed(31'h3f8adc76) * $signed(16'h1);
  assign T6989 = T2943[1'h0:1'h0];
  assign T6990 = T7005 ? twiddle4_3_15_real : twiddle4_3_14_real;
  assign twiddle4_3_14_real = T6996 + T6991;
  assign T6991 = {T6994, T6992};
  assign T6992 = $signed(T6993) / $signed(22'h100000);
  assign T6993 = $signed(29'h8395023) * $signed(16'h0);
  assign T6994 = T6995 ? 2'h3 : 2'h0;
  assign T6995 = T6992[6'h2c:6'h2c];
  assign T6996 = $signed(T6997) / $signed(22'h100000);
  assign T6997 = $signed(31'h3f782c2f) * $signed(16'h1);
  assign twiddle4_3_15_real = T7003 + T6998;
  assign T6998 = {T7001, T6999};
  assign T6999 = $signed(T7000) / $signed(22'h100000);
  assign T7000 = $signed(29'h8cec4a0) * $signed(16'h0);
  assign T7001 = T7002 ? 2'h3 : 2'h0;
  assign T7002 = T6999[6'h2c:6'h2c];
  assign T7003 = $signed(T7004) / $signed(22'h100000);
  assign T7004 = $signed(31'h3f641b8d) * $signed(16'h1);
  assign T7005 = T2943[1'h0:1'h0];
  assign T7006 = T2943[1'h1:1'h1];
  assign T7007 = T2943[2'h2:2'h2];
  assign T7008 = T6938[6'h2e:6'h2e];
  assign T7009 = T2943[2'h3:2'h3];
  assign T7010 = {T7149, T7011};
  assign T7011 = T7148 ? T7082 : T7012;
  assign T7012 = T7081 ? T7047 : T7013;
  assign T7013 = T7046 ? T7030 : T7014;
  assign T7014 = T7029 ? twiddle4_3_17_real : twiddle4_3_16_real;
  assign twiddle4_3_16_real = T7020 + T7015;
  assign T7015 = {T7018, T7016};
  assign T7016 = $signed(T7017) / $signed(22'h100000);
  assign T7017 = $signed(29'h9640837) * $signed(16'h0);
  assign T7018 = T7019 ? 2'h3 : 2'h0;
  assign T7019 = T7016[6'h2c:6'h2c];
  assign T7020 = $signed(T7021) / $signed(22'h100000);
  assign T7021 = $signed(31'h3f4eaafe) * $signed(16'h1);
  assign twiddle4_3_17_real = T7027 + T7022;
  assign T7022 = {T7025, T7023};
  assign T7023 = $signed(T7024) / $signed(22'h100000);
  assign T7024 = $signed(29'h9f917ab) * $signed(16'h0);
  assign T7025 = T7026 ? 2'h3 : 2'h0;
  assign T7026 = T7023[6'h2c:6'h2c];
  assign T7027 = $signed(T7028) / $signed(22'h100000);
  assign T7028 = $signed(31'h3f37daf9) * $signed(16'h1);
  assign T7029 = T2943[1'h0:1'h0];
  assign T7030 = T7045 ? twiddle4_3_19_real : twiddle4_3_18_real;
  assign twiddle4_3_18_real = T7036 + T7031;
  assign T7031 = {T7034, T7032};
  assign T7032 = $signed(T7033) / $signed(22'h100000);
  assign T7033 = $signed(29'ha8defc2) * $signed(16'h0);
  assign T7034 = T7035 ? 2'h3 : 2'h0;
  assign T7035 = T7032[6'h2c:6'h2c];
  assign T7036 = $signed(T7037) / $signed(22'h100000);
  assign T7037 = $signed(31'h3f1fabff) * $signed(16'h1);
  assign twiddle4_3_19_real = T7043 + T7038;
  assign T7038 = {T7041, T7039};
  assign T7039 = $signed(T7040) / $signed(22'h100000);
  assign T7040 = $signed(29'hb228d41) * $signed(16'h0);
  assign T7041 = T7042 ? 2'h3 : 2'h0;
  assign T7042 = T7039[6'h2c:6'h2c];
  assign T7043 = $signed(T7044) / $signed(22'h100000);
  assign T7044 = $signed(31'h3f061e94) * $signed(16'h1);
  assign T7045 = T2943[1'h0:1'h0];
  assign T7046 = T2943[1'h1:1'h1];
  assign T7047 = T7080 ? T7064 : T7048;
  assign T7048 = T7063 ? twiddle4_3_21_real : twiddle4_3_20_real;
  assign twiddle4_3_20_real = T7054 + T7049;
  assign T7049 = {T7052, T7050};
  assign T7050 = $signed(T7051) / $signed(22'h100000);
  assign T7051 = $signed(29'hbb6ecef) * $signed(16'h0);
  assign T7052 = T7053 ? 2'h3 : 2'h0;
  assign T7053 = T7050[6'h2c:6'h2c];
  assign T7054 = $signed(T7055) / $signed(22'h100000);
  assign T7055 = $signed(31'h3eeb3347) * $signed(16'h1);
  assign twiddle4_3_21_real = T7061 + T7056;
  assign T7056 = {T7059, T7057};
  assign T7057 = $signed(T7058) / $signed(22'h100000);
  assign T7058 = $signed(29'hc4b0b93) * $signed(16'h0);
  assign T7059 = T7060 ? 2'h3 : 2'h0;
  assign T7060 = T7057[6'h2c:6'h2c];
  assign T7061 = $signed(T7062) / $signed(22'h100000);
  assign T7062 = $signed(31'h3eceeaad) * $signed(16'h1);
  assign T7063 = T2943[1'h0:1'h0];
  assign T7064 = T7079 ? twiddle4_3_23_real : twiddle4_3_22_real;
  assign twiddle4_3_22_real = T7070 + T7065;
  assign T7065 = {T7068, T7066};
  assign T7066 = $signed(T7067) / $signed(22'h100000);
  assign T7067 = $signed(29'hcdee5f9) * $signed(16'h0);
  assign T7068 = T7069 ? 2'h3 : 2'h0;
  assign T7069 = T7066[6'h2c:6'h2c];
  assign T7070 = $signed(T7071) / $signed(22'h100000);
  assign T7071 = $signed(31'h3eb14562) * $signed(16'h1);
  assign twiddle4_3_23_real = T7077 + T7072;
  assign T7072 = {T7075, T7073};
  assign T7073 = $signed(T7074) / $signed(22'h100000);
  assign T7074 = $signed(29'hd7278ea) * $signed(16'h0);
  assign T7075 = T7076 ? 2'h3 : 2'h0;
  assign T7076 = T7073[6'h2c:6'h2c];
  assign T7077 = $signed(T7078) / $signed(22'h100000);
  assign T7078 = $signed(31'h3e92440d) * $signed(16'h1);
  assign T7079 = T2943[1'h0:1'h0];
  assign T7080 = T2943[1'h1:1'h1];
  assign T7081 = T2943[2'h2:2'h2];
  assign T7082 = T7147 ? T7117 : T7083;
  assign T7083 = T7116 ? T7100 : T7084;
  assign T7084 = T7099 ? twiddle4_3_25_real : twiddle4_3_24_real;
  assign twiddle4_3_24_real = T7090 + T7085;
  assign T7085 = {T7088, T7086};
  assign T7086 = $signed(T7087) / $signed(22'h100000);
  assign T7087 = $signed(29'he05c135) * $signed(16'h0);
  assign T7088 = T7089 ? 2'h3 : 2'h0;
  assign T7089 = T7086[6'h2c:6'h2c];
  assign T7090 = $signed(T7091) / $signed(22'h100000);
  assign T7091 = $signed(31'h3e71e758) * $signed(16'h1);
  assign twiddle4_3_25_real = T7097 + T7092;
  assign T7092 = {T7095, T7093};
  assign T7093 = $signed(T7094) / $signed(22'h100000);
  assign T7094 = $signed(29'he98bba6) * $signed(16'h0);
  assign T7095 = T7096 ? 2'h3 : 2'h0;
  assign T7096 = T7093[6'h2c:6'h2c];
  assign T7097 = $signed(T7098) / $signed(22'h100000);
  assign T7098 = $signed(31'h3e502ff8) * $signed(16'h1);
  assign T7099 = T2943[1'h0:1'h0];
  assign T7100 = T7115 ? twiddle4_3_27_real : twiddle4_3_26_real;
  assign twiddle4_3_26_real = T7106 + T7101;
  assign T7101 = {T7104, T7102};
  assign T7102 = $signed(T7103) / $signed(22'h100000);
  assign T7103 = $signed(29'hf2b650f) * $signed(16'h0);
  assign T7104 = T7105 ? 2'h3 : 2'h0;
  assign T7105 = T7102[6'h2c:6'h2c];
  assign T7106 = $signed(T7107) / $signed(22'h100000);
  assign T7107 = $signed(31'h3e2d1ea7) * $signed(16'h1);
  assign twiddle4_3_27_real = T7113 + T7108;
  assign T7108 = {T7111, T7109};
  assign T7109 = $signed(T7110) / $signed(22'h100000);
  assign T7110 = $signed(29'hfbdba40) * $signed(16'h0);
  assign T7111 = T7112 ? 2'h3 : 2'h0;
  assign T7112 = T7109[6'h2c:6'h2c];
  assign T7113 = $signed(T7114) / $signed(22'h100000);
  assign T7114 = $signed(31'h3e08b429) * $signed(16'h1);
  assign T7115 = T2943[1'h0:1'h0];
  assign T7116 = T2943[1'h1:1'h1];
  assign T7117 = T7146 ? T7132 : T7118;
  assign T7118 = T7131 ? twiddle4_3_29_real : twiddle4_3_28_real;
  assign twiddle4_3_28_real = T7123 + T7119;
  assign T7119 = {T7122, T7120};
  assign T7120 = $signed(T7121) / $signed(22'h100000);
  assign T7121 = $signed(30'h104fb80e) * $signed(16'h0);
  assign T7122 = T7120[6'h2d:6'h2d];
  assign T7123 = $signed(T7124) / $signed(22'h100000);
  assign T7124 = $signed(31'h3de2f147) * $signed(16'h1);
  assign twiddle4_3_29_real = T7129 + T7125;
  assign T7125 = {T7128, T7126};
  assign T7126 = $signed(T7127) / $signed(22'h100000);
  assign T7127 = $signed(30'h10e15b4e) * $signed(16'h0);
  assign T7128 = T7126[6'h2d:6'h2d];
  assign T7129 = $signed(T7130) / $signed(22'h100000);
  assign T7130 = $signed(31'h3dbbd6d4) * $signed(16'h1);
  assign T7131 = T2943[1'h0:1'h0];
  assign T7132 = T7145 ? twiddle4_3_31_real : twiddle4_3_30_real;
  assign twiddle4_3_30_real = T7137 + T7133;
  assign T7133 = {T7136, T7134};
  assign T7134 = $signed(T7135) / $signed(22'h100000);
  assign T7135 = $signed(30'h1172a0d7) * $signed(16'h0);
  assign T7136 = T7134[6'h2d:6'h2d];
  assign T7137 = $signed(T7138) / $signed(22'h100000);
  assign T7138 = $signed(31'h3d9365a7) * $signed(16'h1);
  assign twiddle4_3_31_real = T7143 + T7139;
  assign T7139 = {T7142, T7140};
  assign T7140 = $signed(T7141) / $signed(22'h100000);
  assign T7141 = $signed(30'h12038583) * $signed(16'h0);
  assign T7142 = T7140[6'h2d:6'h2d];
  assign T7143 = $signed(T7144) / $signed(22'h100000);
  assign T7144 = $signed(31'h3d699ea2) * $signed(16'h1);
  assign T7145 = T2943[1'h0:1'h0];
  assign T7146 = T2943[1'h1:1'h1];
  assign T7147 = T2943[2'h2:2'h2];
  assign T7148 = T2943[2'h3:2'h3];
  assign T7149 = T7011[6'h2e:6'h2e];
  assign T7150 = T2943[3'h4:3'h4];
  assign T7151 = {T7392, T7152};
  assign T7152 = T7391 ? T7279 : T7153;
  assign T7153 = T7278 ? T7216 : T7154;
  assign T7154 = T7215 ? T7185 : T7155;
  assign T7155 = T7184 ? T7170 : T7156;
  assign T7156 = T7169 ? twiddle4_3_33_real : twiddle4_3_32_real;
  assign twiddle4_3_32_real = T7161 + T7157;
  assign T7157 = {T7160, T7158};
  assign T7158 = $signed(T7159) / $signed(22'h100000);
  assign T7159 = $signed(30'h1294062e) * $signed(16'h0);
  assign T7160 = T7158[6'h2d:6'h2d];
  assign T7161 = $signed(T7162) / $signed(22'h100000);
  assign T7162 = $signed(31'h3d3e82ad) * $signed(16'h1);
  assign twiddle4_3_33_real = T7167 + T7163;
  assign T7163 = {T7166, T7164};
  assign T7164 = $signed(T7165) / $signed(22'h100000);
  assign T7165 = $signed(30'h13241fb6) * $signed(16'h0);
  assign T7166 = T7164[6'h2d:6'h2d];
  assign T7167 = $signed(T7168) / $signed(22'h100000);
  assign T7168 = $signed(31'h3d1212b7) * $signed(16'h1);
  assign T7169 = T2943[1'h0:1'h0];
  assign T7170 = T7183 ? twiddle4_3_35_real : twiddle4_3_34_real;
  assign twiddle4_3_34_real = T7175 + T7171;
  assign T7171 = {T7174, T7172};
  assign T7172 = $signed(T7173) / $signed(22'h100000);
  assign T7173 = $signed(30'h13b3cefa) * $signed(16'h0);
  assign T7174 = T7172[6'h2d:6'h2d];
  assign T7175 = $signed(T7176) / $signed(22'h100000);
  assign T7176 = $signed(31'h3ce44fb6) * $signed(16'h1);
  assign twiddle4_3_35_real = T7181 + T7177;
  assign T7177 = {T7180, T7178};
  assign T7178 = $signed(T7179) / $signed(22'h100000);
  assign T7179 = $signed(30'h144310dc) * $signed(16'h0);
  assign T7180 = T7178[6'h2d:6'h2d];
  assign T7181 = $signed(T7182) / $signed(22'h100000);
  assign T7182 = $signed(31'h3cb53aaa) * $signed(16'h1);
  assign T7183 = T2943[1'h0:1'h0];
  assign T7184 = T2943[1'h1:1'h1];
  assign T7185 = T7214 ? T7200 : T7186;
  assign T7186 = T7199 ? twiddle4_3_37_real : twiddle4_3_36_real;
  assign twiddle4_3_36_real = T7191 + T7187;
  assign T7187 = {T7190, T7188};
  assign T7188 = $signed(T7189) / $signed(22'h100000);
  assign T7189 = $signed(30'h14d1e242) * $signed(16'h0);
  assign T7190 = T7188[6'h2d:6'h2d];
  assign T7191 = $signed(T7192) / $signed(22'h100000);
  assign T7192 = $signed(31'h3c84d496) * $signed(16'h1);
  assign twiddle4_3_37_real = T7197 + T7193;
  assign T7193 = {T7196, T7194};
  assign T7194 = $signed(T7195) / $signed(22'h100000);
  assign T7195 = $signed(30'h15604012) * $signed(16'h0);
  assign T7196 = T7194[6'h2d:6'h2d];
  assign T7197 = $signed(T7198) / $signed(22'h100000);
  assign T7198 = $signed(31'h3c531e88) * $signed(16'h1);
  assign T7199 = T2943[1'h0:1'h0];
  assign T7200 = T7213 ? twiddle4_3_39_real : twiddle4_3_38_real;
  assign twiddle4_3_38_real = T7205 + T7201;
  assign T7201 = {T7204, T7202};
  assign T7202 = $signed(T7203) / $signed(22'h100000);
  assign T7203 = $signed(30'h15ee2737) * $signed(16'h0);
  assign T7204 = T7202[6'h2d:6'h2d];
  assign T7205 = $signed(T7206) / $signed(22'h100000);
  assign T7206 = $signed(31'h3c201994) * $signed(16'h1);
  assign twiddle4_3_39_real = T7211 + T7207;
  assign T7207 = {T7210, T7208};
  assign T7208 = $signed(T7209) / $signed(22'h100000);
  assign T7209 = $signed(30'h167b949c) * $signed(16'h0);
  assign T7210 = T7208[6'h2d:6'h2d];
  assign T7211 = $signed(T7212) / $signed(22'h100000);
  assign T7212 = $signed(31'h3bebc6d5) * $signed(16'h1);
  assign T7213 = T2943[1'h0:1'h0];
  assign T7214 = T2943[1'h1:1'h1];
  assign T7215 = T2943[2'h2:2'h2];
  assign T7216 = T7277 ? T7247 : T7217;
  assign T7217 = T7246 ? T7232 : T7218;
  assign T7218 = T7231 ? twiddle4_3_41_real : twiddle4_3_40_real;
  assign twiddle4_3_40_real = T7223 + T7219;
  assign T7219 = {T7222, T7220};
  assign T7220 = $signed(T7221) / $signed(22'h100000);
  assign T7221 = $signed(30'h17088530) * $signed(16'h0);
  assign T7222 = T7220[6'h2d:6'h2d];
  assign T7223 = $signed(T7224) / $signed(22'h100000);
  assign T7224 = $signed(31'h3bb6276d) * $signed(16'h1);
  assign twiddle4_3_41_real = T7229 + T7225;
  assign T7225 = {T7228, T7226};
  assign T7226 = $signed(T7227) / $signed(22'h100000);
  assign T7227 = $signed(30'h1794f5e6) * $signed(16'h0);
  assign T7228 = T7226[6'h2d:6'h2d];
  assign T7229 = $signed(T7230) / $signed(22'h100000);
  assign T7230 = $signed(31'h3b7f3c87) * $signed(16'h1);
  assign T7231 = T2943[1'h0:1'h0];
  assign T7232 = T7245 ? twiddle4_3_43_real : twiddle4_3_42_real;
  assign twiddle4_3_42_real = T7237 + T7233;
  assign T7233 = {T7236, T7234};
  assign T7234 = $signed(T7235) / $signed(22'h100000);
  assign T7235 = $signed(30'h1820e3b0) * $signed(16'h0);
  assign T7236 = T7234[6'h2d:6'h2d];
  assign T7237 = $signed(T7238) / $signed(22'h100000);
  assign T7238 = $signed(31'h3b470752) * $signed(16'h1);
  assign twiddle4_3_43_real = T7243 + T7239;
  assign T7239 = {T7242, T7240};
  assign T7240 = $signed(T7241) / $signed(22'h100000);
  assign T7241 = $signed(30'h18ac4b86) * $signed(16'h0);
  assign T7242 = T7240[6'h2d:6'h2d];
  assign T7243 = $signed(T7244) / $signed(22'h100000);
  assign T7244 = $signed(31'h3b0d8908) * $signed(16'h1);
  assign T7245 = T2943[1'h0:1'h0];
  assign T7246 = T2943[1'h1:1'h1];
  assign T7247 = T7276 ? T7262 : T7248;
  assign T7248 = T7261 ? twiddle4_3_45_real : twiddle4_3_44_real;
  assign twiddle4_3_44_real = T7253 + T7249;
  assign T7249 = {T7252, T7250};
  assign T7250 = $signed(T7251) / $signed(22'h100000);
  assign T7251 = $signed(30'h19372a63) * $signed(16'h0);
  assign T7252 = T7250[6'h2d:6'h2d];
  assign T7253 = $signed(T7254) / $signed(22'h100000);
  assign T7254 = $signed(31'h3ad2c2e7) * $signed(16'h1);
  assign twiddle4_3_45_real = T7259 + T7255;
  assign T7255 = {T7258, T7256};
  assign T7256 = $signed(T7257) / $signed(22'h100000);
  assign T7257 = $signed(30'h19c17d44) * $signed(16'h0);
  assign T7258 = T7256[6'h2d:6'h2d];
  assign T7259 = $signed(T7260) / $signed(22'h100000);
  assign T7260 = $signed(31'h3a96b636) * $signed(16'h1);
  assign T7261 = T2943[1'h0:1'h0];
  assign T7262 = T7275 ? twiddle4_3_47_real : twiddle4_3_46_real;
  assign twiddle4_3_46_real = T7267 + T7263;
  assign T7263 = {T7266, T7264};
  assign T7264 = $signed(T7265) / $signed(22'h100000);
  assign T7265 = $signed(30'h1a4b4127) * $signed(16'h0);
  assign T7266 = T7264[6'h2d:6'h2d];
  assign T7267 = $signed(T7268) / $signed(22'h100000);
  assign T7268 = $signed(31'h3a596441) * $signed(16'h1);
  assign twiddle4_3_47_real = T7273 + T7269;
  assign T7269 = {T7272, T7270};
  assign T7270 = $signed(T7271) / $signed(22'h100000);
  assign T7271 = $signed(30'h1ad47312) * $signed(16'h0);
  assign T7272 = T7270[6'h2d:6'h2d];
  assign T7273 = $signed(T7274) / $signed(22'h100000);
  assign T7274 = $signed(31'h3a1ace5e) * $signed(16'h1);
  assign T7275 = T2943[1'h0:1'h0];
  assign T7276 = T2943[1'h1:1'h1];
  assign T7277 = T2943[2'h2:2'h2];
  assign T7278 = T2943[2'h3:2'h3];
  assign T7279 = T7390 ? T7342 : T7280;
  assign T7280 = T7341 ? T7311 : T7281;
  assign T7281 = T7310 ? T7296 : T7282;
  assign T7282 = T7295 ? twiddle4_3_49_real : twiddle4_3_48_real;
  assign twiddle4_3_48_real = T7287 + T7283;
  assign T7283 = {T7286, T7284};
  assign T7284 = $signed(T7285) / $signed(22'h100000);
  assign T7285 = $signed(30'h1b5d1009) * $signed(16'h0);
  assign T7286 = T7284[6'h2d:6'h2d];
  assign T7287 = $signed(T7288) / $signed(22'h100000);
  assign T7288 = $signed(31'h39daf5e8) * $signed(16'h1);
  assign twiddle4_3_49_real = T7293 + T7289;
  assign T7289 = {T7292, T7290};
  assign T7290 = $signed(T7291) / $signed(22'h100000);
  assign T7291 = $signed(30'h1be51517) * $signed(16'h0);
  assign T7292 = T7290[6'h2d:6'h2d];
  assign T7293 = $signed(T7294) / $signed(22'h100000);
  assign T7294 = $signed(31'h3999dc41) * $signed(16'h1);
  assign T7295 = T2943[1'h0:1'h0];
  assign T7296 = T7309 ? twiddle4_3_51_real : twiddle4_3_50_real;
  assign twiddle4_3_50_real = T7301 + T7297;
  assign T7297 = {T7300, T7298};
  assign T7298 = $signed(T7299) / $signed(22'h100000);
  assign T7299 = $signed(30'h1c6c7f49) * $signed(16'h0);
  assign T7300 = T7298[6'h2d:6'h2d];
  assign T7301 = $signed(T7302) / $signed(22'h100000);
  assign T7302 = $signed(31'h395782d3) * $signed(16'h1);
  assign twiddle4_3_51_real = T7307 + T7303;
  assign T7303 = {T7306, T7304};
  assign T7304 = $signed(T7305) / $signed(22'h100000);
  assign T7305 = $signed(30'h1cf34bae) * $signed(16'h0);
  assign T7306 = T7304[6'h2d:6'h2d];
  assign T7307 = $signed(T7308) / $signed(22'h100000);
  assign T7308 = $signed(31'h3913eb0e) * $signed(16'h1);
  assign T7309 = T2943[1'h0:1'h0];
  assign T7310 = T2943[1'h1:1'h1];
  assign T7311 = T7340 ? T7326 : T7312;
  assign T7312 = T7325 ? twiddle4_3_53_real : twiddle4_3_52_real;
  assign twiddle4_3_52_real = T7317 + T7313;
  assign T7313 = {T7316, T7314};
  assign T7314 = $signed(T7315) / $signed(22'h100000);
  assign T7315 = $signed(30'h1d79775b) * $signed(16'h0);
  assign T7316 = T7314[6'h2d:6'h2d];
  assign T7317 = $signed(T7318) / $signed(22'h100000);
  assign T7318 = $signed(31'h38cf1669) * $signed(16'h1);
  assign twiddle4_3_53_real = T7323 + T7319;
  assign T7319 = {T7322, T7320};
  assign T7320 = $signed(T7321) / $signed(22'h100000);
  assign T7321 = $signed(30'h1dfeff66) * $signed(16'h0);
  assign T7322 = T7320[6'h2d:6'h2d];
  assign T7323 = $signed(T7324) / $signed(22'h100000);
  assign T7324 = $signed(31'h38890662) * $signed(16'h1);
  assign T7325 = T2943[1'h0:1'h0];
  assign T7326 = T7339 ? twiddle4_3_55_real : twiddle4_3_54_real;
  assign twiddle4_3_54_real = T7331 + T7327;
  assign T7327 = {T7330, T7328};
  assign T7328 = $signed(T7329) / $signed(22'h100000);
  assign T7329 = $signed(30'h1e83e0ea) * $signed(16'h0);
  assign T7330 = T7328[6'h2d:6'h2d];
  assign T7331 = $signed(T7332) / $signed(22'h100000);
  assign T7332 = $signed(31'h3841bc7f) * $signed(16'h1);
  assign twiddle4_3_55_real = T7337 + T7333;
  assign T7333 = {T7336, T7334};
  assign T7334 = $signed(T7335) / $signed(22'h100000);
  assign T7335 = $signed(30'h1f081906) * $signed(16'h0);
  assign T7336 = T7334[6'h2d:6'h2d];
  assign T7337 = $signed(T7338) / $signed(22'h100000);
  assign T7338 = $signed(31'h37f93a4b) * $signed(16'h1);
  assign T7339 = T2943[1'h0:1'h0];
  assign T7340 = T2943[1'h1:1'h1];
  assign T7341 = T2943[2'h2:2'h2];
  assign T7342 = T7389 ? T7367 : T7343;
  assign T7343 = T7366 ? T7356 : T7344;
  assign T7344 = T7355 ? twiddle4_3_57_real : twiddle4_3_56_real;
  assign twiddle4_3_56_real = T7349 + T7345;
  assign T7345 = {T7348, T7346};
  assign T7346 = $signed(T7347) / $signed(22'h100000);
  assign T7347 = $signed(30'h1f8ba4db) * $signed(16'h0);
  assign T7348 = T7346[6'h2d:6'h2d];
  assign T7349 = $signed(T7350) / $signed(22'h100000);
  assign T7350 = $signed(31'h37af8158) * $signed(16'h1);
  assign twiddle4_3_57_real = T7353 + T7351;
  assign T7351 = $signed(T7352) / $signed(22'h100000);
  assign T7352 = $signed(31'h200e8190) * $signed(16'h0);
  assign T7353 = $signed(T7354) / $signed(22'h100000);
  assign T7354 = $signed(31'h37649341) * $signed(16'h1);
  assign T7355 = T2943[1'h0:1'h0];
  assign T7356 = T7365 ? twiddle4_3_59_real : twiddle4_3_58_real;
  assign twiddle4_3_58_real = T7359 + T7357;
  assign T7357 = $signed(T7358) / $signed(22'h100000);
  assign T7358 = $signed(31'h2090ac4d) * $signed(16'h0);
  assign T7359 = $signed(T7360) / $signed(22'h100000);
  assign T7360 = $signed(31'h371871a4) * $signed(16'h1);
  assign twiddle4_3_59_real = T7363 + T7361;
  assign T7361 = $signed(T7362) / $signed(22'h100000);
  assign T7362 = $signed(31'h21122240) * $signed(16'h0);
  assign T7363 = $signed(T7364) / $signed(22'h100000);
  assign T7364 = $signed(31'h36cb1e29) * $signed(16'h1);
  assign T7365 = T2943[1'h0:1'h0];
  assign T7366 = T2943[1'h1:1'h1];
  assign T7367 = T7388 ? T7378 : T7368;
  assign T7368 = T7377 ? twiddle4_3_61_real : twiddle4_3_60_real;
  assign twiddle4_3_60_real = T7371 + T7369;
  assign T7369 = $signed(T7370) / $signed(22'h100000);
  assign T7370 = $signed(31'h2192e09a) * $signed(16'h0);
  assign T7371 = $signed(T7372) / $signed(22'h100000);
  assign T7372 = $signed(31'h367c9a7d) * $signed(16'h1);
  assign twiddle4_3_61_real = T7375 + T7373;
  assign T7373 = $signed(T7374) / $signed(22'h100000);
  assign T7374 = $signed(31'h2212e491) * $signed(16'h0);
  assign T7375 = $signed(T7376) / $signed(22'h100000);
  assign T7376 = $signed(31'h362ce854) * $signed(16'h1);
  assign T7377 = T2943[1'h0:1'h0];
  assign T7378 = T7387 ? twiddle4_3_63_real : twiddle4_3_62_real;
  assign twiddle4_3_62_real = T7381 + T7379;
  assign T7379 = $signed(T7380) / $signed(22'h100000);
  assign T7380 = $signed(31'h22922b5e) * $signed(16'h0);
  assign T7381 = $signed(T7382) / $signed(22'h100000);
  assign T7382 = $signed(31'h35dc0968) * $signed(16'h1);
  assign twiddle4_3_63_real = T7385 + T7383;
  assign T7383 = $signed(T7384) / $signed(22'h100000);
  assign T7384 = $signed(31'h2310b23e) * $signed(16'h0);
  assign T7385 = $signed(T7386) / $signed(22'h100000);
  assign T7386 = $signed(31'h3589ff7a) * $signed(16'h1);
  assign T7387 = T2943[1'h0:1'h0];
  assign T7388 = T2943[1'h1:1'h1];
  assign T7389 = T2943[2'h2:2'h2];
  assign T7390 = T2943[2'h3:2'h3];
  assign T7391 = T2943[3'h4:3'h4];
  assign T7392 = T7152[6'h2e:6'h2e];
  assign T7393 = T2943[3'h5:3'h5];
  assign T7394 = {T7805, T7395};
  assign T7395 = T7804 ? T7586 : T7396;
  assign T7396 = T7585 ? T7491 : T7397;
  assign T7397 = T7490 ? T7444 : T7398;
  assign T7398 = T7443 ? T7421 : T7399;
  assign T7399 = T7420 ? T7410 : T7400;
  assign T7400 = T7409 ? twiddle4_3_65_real : twiddle4_3_64_real;
  assign twiddle4_3_64_real = T7403 + T7401;
  assign T7401 = $signed(T7402) / $signed(22'h100000);
  assign T7402 = $signed(31'h238e7673) * $signed(16'h0);
  assign T7403 = $signed(T7404) / $signed(22'h100000);
  assign T7404 = $signed(31'h3536cc52) * $signed(16'h1);
  assign twiddle4_3_65_real = T7407 + T7405;
  assign T7405 = $signed(T7406) / $signed(22'h100000);
  assign T7406 = $signed(31'h240b7542) * $signed(16'h0);
  assign T7407 = $signed(T7408) / $signed(22'h100000);
  assign T7408 = $signed(31'h34e271bd) * $signed(16'h1);
  assign T7409 = T2943[1'h0:1'h0];
  assign T7410 = T7419 ? twiddle4_3_67_real : twiddle4_3_66_real;
  assign twiddle4_3_66_real = T7413 + T7411;
  assign T7411 = $signed(T7412) / $signed(22'h100000);
  assign T7412 = $signed(31'h2487abf7) * $signed(16'h0);
  assign T7413 = $signed(T7414) / $signed(22'h100000);
  assign T7414 = $signed(31'h348cf190) * $signed(16'h1);
  assign twiddle4_3_67_real = T7417 + T7415;
  assign T7415 = $signed(T7416) / $signed(22'h100000);
  assign T7416 = $signed(31'h250317de) * $signed(16'h0);
  assign T7417 = $signed(T7418) / $signed(22'h100000);
  assign T7418 = $signed(31'h34364da5) * $signed(16'h1);
  assign T7419 = T2943[1'h0:1'h0];
  assign T7420 = T2943[1'h1:1'h1];
  assign T7421 = T7442 ? T7432 : T7422;
  assign T7422 = T7431 ? twiddle4_3_69_real : twiddle4_3_68_real;
  assign twiddle4_3_68_real = T7425 + T7423;
  assign T7423 = $signed(T7424) / $signed(22'h100000);
  assign T7424 = $signed(31'h257db64b) * $signed(16'h0);
  assign T7425 = $signed(T7426) / $signed(22'h100000);
  assign T7426 = $signed(31'h33de87de) * $signed(16'h1);
  assign twiddle4_3_69_real = T7429 + T7427;
  assign T7427 = $signed(T7428) / $signed(22'h100000);
  assign T7428 = $signed(31'h25f78496) * $signed(16'h0);
  assign T7429 = $signed(T7430) / $signed(22'h100000);
  assign T7430 = $signed(31'h3385a221) * $signed(16'h1);
  assign T7431 = T2943[1'h0:1'h0];
  assign T7432 = T7441 ? twiddle4_3_71_real : twiddle4_3_70_real;
  assign twiddle4_3_70_real = T7435 + T7433;
  assign T7433 = $signed(T7434) / $signed(22'h100000);
  assign T7434 = $signed(31'h2670801a) * $signed(16'h0);
  assign T7435 = $signed(T7436) / $signed(22'h100000);
  assign T7436 = $signed(31'h332b9e5d) * $signed(16'h1);
  assign twiddle4_3_71_real = T7439 + T7437;
  assign T7437 = $signed(T7438) / $signed(22'h100000);
  assign T7438 = $signed(31'h26e8a637) * $signed(16'h0);
  assign T7439 = $signed(T7440) / $signed(22'h100000);
  assign T7440 = $signed(31'h32d07e85) * $signed(16'h1);
  assign T7441 = T2943[1'h0:1'h0];
  assign T7442 = T2943[1'h1:1'h1];
  assign T7443 = T2943[2'h2:2'h2];
  assign T7444 = T7489 ? T7467 : T7445;
  assign T7445 = T7466 ? T7456 : T7446;
  assign T7446 = T7455 ? twiddle4_3_73_real : twiddle4_3_72_real;
  assign twiddle4_3_72_real = T7449 + T7447;
  assign T7447 = $signed(T7448) / $signed(22'h100000);
  assign T7448 = $signed(31'h275ff452) * $signed(16'h0);
  assign T7449 = $signed(T7450) / $signed(22'h100000);
  assign T7450 = $signed(31'h32744493) * $signed(16'h1);
  assign twiddle4_3_73_real = T7453 + T7451;
  assign T7451 = $signed(T7452) / $signed(22'h100000);
  assign T7452 = $signed(31'h27d667d5) * $signed(16'h0);
  assign T7453 = $signed(T7454) / $signed(22'h100000);
  assign T7454 = $signed(31'h3216f286) * $signed(16'h1);
  assign T7455 = T2943[1'h0:1'h0];
  assign T7456 = T7465 ? twiddle4_3_75_real : twiddle4_3_74_real;
  assign twiddle4_3_74_real = T7459 + T7457;
  assign T7457 = $signed(T7458) / $signed(22'h100000);
  assign T7458 = $signed(31'h284bfe2f) * $signed(16'h0);
  assign T7459 = $signed(T7460) / $signed(22'h100000);
  assign T7460 = $signed(31'h31b88a66) * $signed(16'h1);
  assign twiddle4_3_75_real = T7463 + T7461;
  assign T7461 = $signed(T7462) / $signed(22'h100000);
  assign T7462 = $signed(31'h28c0b4d2) * $signed(16'h0);
  assign T7463 = $signed(T7464) / $signed(22'h100000);
  assign T7464 = $signed(31'h31590e3d) * $signed(16'h1);
  assign T7465 = T2943[1'h0:1'h0];
  assign T7466 = T2943[1'h1:1'h1];
  assign T7467 = T7488 ? T7478 : T7468;
  assign T7468 = T7477 ? twiddle4_3_77_real : twiddle4_3_76_real;
  assign twiddle4_3_76_real = T7471 + T7469;
  assign T7469 = $signed(T7470) / $signed(22'h100000);
  assign T7470 = $signed(31'h29348937) * $signed(16'h0);
  assign T7471 = $signed(T7472) / $signed(22'h100000);
  assign T7472 = $signed(31'h30f8801f) * $signed(16'h1);
  assign twiddle4_3_77_real = T7475 + T7473;
  assign T7473 = $signed(T7474) / $signed(22'h100000);
  assign T7474 = $signed(31'h29a778da) * $signed(16'h0);
  assign T7475 = $signed(T7476) / $signed(22'h100000);
  assign T7476 = $signed(31'h3096e223) * $signed(16'h1);
  assign T7477 = T2943[1'h0:1'h0];
  assign T7478 = T7487 ? twiddle4_3_79_real : twiddle4_3_78_real;
  assign twiddle4_3_78_real = T7481 + T7479;
  assign T7479 = $signed(T7480) / $signed(22'h100000);
  assign T7480 = $signed(31'h2a19813e) * $signed(16'h0);
  assign T7481 = $signed(T7482) / $signed(22'h100000);
  assign T7482 = $signed(31'h30343667) * $signed(16'h1);
  assign twiddle4_3_79_real = T7485 + T7483;
  assign T7483 = $signed(T7484) / $signed(22'h100000);
  assign T7484 = $signed(31'h2a8a9fea) * $signed(16'h0);
  assign T7485 = $signed(T7486) / $signed(22'h100000);
  assign T7486 = $signed(31'h2fd07f0f) * $signed(16'h1);
  assign T7487 = T2943[1'h0:1'h0];
  assign T7488 = T2943[1'h1:1'h1];
  assign T7489 = T2943[2'h2:2'h2];
  assign T7490 = T2943[2'h3:2'h3];
  assign T7491 = T7584 ? T7538 : T7492;
  assign T7492 = T7537 ? T7515 : T7493;
  assign T7493 = T7514 ? T7504 : T7494;
  assign T7494 = T7503 ? twiddle4_3_81_real : twiddle4_3_80_real;
  assign twiddle4_3_80_real = T7497 + T7495;
  assign T7495 = $signed(T7496) / $signed(22'h100000);
  assign T7496 = $signed(31'h2afad269) * $signed(16'h0);
  assign T7497 = $signed(T7498) / $signed(22'h100000);
  assign T7498 = $signed(31'h2f6bbe44) * $signed(16'h1);
  assign twiddle4_3_81_real = T7501 + T7499;
  assign T7499 = $signed(T7500) / $signed(22'h100000);
  assign T7500 = $signed(31'h2b6a164c) * $signed(16'h0);
  assign T7501 = $signed(T7502) / $signed(22'h100000);
  assign T7502 = $signed(31'h2f05f637) * $signed(16'h1);
  assign T7503 = T2943[1'h0:1'h0];
  assign T7504 = T7513 ? twiddle4_3_83_real : twiddle4_3_82_real;
  assign twiddle4_3_82_real = T7507 + T7505;
  assign T7505 = $signed(T7506) / $signed(22'h100000);
  assign T7506 = $signed(31'h2bd8692b) * $signed(16'h0);
  assign T7507 = $signed(T7508) / $signed(22'h100000);
  assign T7508 = $signed(31'h2e9f291b) * $signed(16'h1);
  assign twiddle4_3_83_real = T7511 + T7509;
  assign T7509 = $signed(T7510) / $signed(22'h100000);
  assign T7510 = $signed(31'h2c45c89f) * $signed(16'h0);
  assign T7511 = $signed(T7512) / $signed(22'h100000);
  assign T7512 = $signed(31'h2e37592c) * $signed(16'h1);
  assign T7513 = T2943[1'h0:1'h0];
  assign T7514 = T2943[1'h1:1'h1];
  assign T7515 = T7536 ? T7526 : T7516;
  assign T7516 = T7525 ? twiddle4_3_85_real : twiddle4_3_84_real;
  assign twiddle4_3_84_real = T7519 + T7517;
  assign T7517 = $signed(T7518) / $signed(22'h100000);
  assign T7518 = $signed(31'h2cb2324b) * $signed(16'h0);
  assign T7519 = $signed(T7520) / $signed(22'h100000);
  assign T7520 = $signed(31'h2dce88a9) * $signed(16'h1);
  assign twiddle4_3_85_real = T7523 + T7521;
  assign T7521 = $signed(T7522) / $signed(22'h100000);
  assign T7522 = $signed(31'h2d1da3d5) * $signed(16'h0);
  assign T7523 = $signed(T7524) / $signed(22'h100000);
  assign T7524 = $signed(31'h2d64b9da) * $signed(16'h1);
  assign T7525 = T2943[1'h0:1'h0];
  assign T7526 = T7535 ? twiddle4_3_87_real : twiddle4_3_86_real;
  assign twiddle4_3_86_real = T7529 + T7527;
  assign T7527 = $signed(T7528) / $signed(22'h100000);
  assign T7528 = $signed(31'h2d881ae7) * $signed(16'h0);
  assign T7529 = $signed(T7530) / $signed(22'h100000);
  assign T7530 = $signed(31'h2cf9ef09) * $signed(16'h1);
  assign twiddle4_3_87_real = T7533 + T7531;
  assign T7531 = $signed(T7532) / $signed(22'h100000);
  assign T7532 = $signed(31'h2df19533) * $signed(16'h0);
  assign T7533 = $signed(T7534) / $signed(22'h100000);
  assign T7534 = $signed(31'h2c8e2a86) * $signed(16'h1);
  assign T7535 = T2943[1'h0:1'h0];
  assign T7536 = T2943[1'h1:1'h1];
  assign T7537 = T2943[2'h2:2'h2];
  assign T7538 = T7583 ? T7561 : T7539;
  assign T7539 = T7560 ? T7550 : T7540;
  assign T7540 = T7549 ? twiddle4_3_89_real : twiddle4_3_88_real;
  assign twiddle4_3_88_real = T7543 + T7541;
  assign T7541 = $signed(T7542) / $signed(22'h100000);
  assign T7542 = $signed(31'h2e5a106f) * $signed(16'h0);
  assign T7543 = $signed(T7544) / $signed(22'h100000);
  assign T7544 = $signed(31'h2c216eaa) * $signed(16'h1);
  assign twiddle4_3_89_real = T7547 + T7545;
  assign T7545 = $signed(T7546) / $signed(22'h100000);
  assign T7546 = $signed(31'h2ec18a58) * $signed(16'h0);
  assign T7547 = $signed(T7548) / $signed(22'h100000);
  assign T7548 = $signed(31'h2bb3bdce) * $signed(16'h1);
  assign T7549 = T2943[1'h0:1'h0];
  assign T7550 = T7559 ? twiddle4_3_91_real : twiddle4_3_90_real;
  assign twiddle4_3_90_real = T7553 + T7551;
  assign T7551 = $signed(T7552) / $signed(22'h100000);
  assign T7552 = $signed(31'h2f2800ae) * $signed(16'h0);
  assign T7553 = $signed(T7554) / $signed(22'h100000);
  assign T7554 = $signed(31'h2b451a54) * $signed(16'h1);
  assign twiddle4_3_91_real = T7557 + T7555;
  assign T7555 = $signed(T7556) / $signed(22'h100000);
  assign T7556 = $signed(31'h2f8d7139) * $signed(16'h0);
  assign T7557 = $signed(T7558) / $signed(22'h100000);
  assign T7558 = $signed(31'h2ad586a3) * $signed(16'h1);
  assign T7559 = T2943[1'h0:1'h0];
  assign T7560 = T2943[1'h1:1'h1];
  assign T7561 = T7582 ? T7572 : T7562;
  assign T7562 = T7571 ? twiddle4_3_93_real : twiddle4_3_92_real;
  assign twiddle4_3_92_real = T7565 + T7563;
  assign T7563 = $signed(T7564) / $signed(22'h100000);
  assign T7564 = $signed(31'h2ff1d9c6) * $signed(16'h0);
  assign T7565 = $signed(T7566) / $signed(22'h100000);
  assign T7566 = $signed(31'h2a650525) * $signed(16'h1);
  assign twiddle4_3_93_real = T7569 + T7567;
  assign T7567 = $signed(T7568) / $signed(22'h100000);
  assign T7568 = $signed(31'h30553827) * $signed(16'h0);
  assign T7569 = $signed(T7570) / $signed(22'h100000);
  assign T7570 = $signed(31'h29f3984b) * $signed(16'h1);
  assign T7571 = T2943[1'h0:1'h0];
  assign T7572 = T7581 ? twiddle4_3_95_real : twiddle4_3_94_real;
  assign twiddle4_3_94_real = T7575 + T7573;
  assign T7573 = $signed(T7574) / $signed(22'h100000);
  assign T7574 = $signed(31'h30b78a35) * $signed(16'h0);
  assign T7575 = $signed(T7576) / $signed(22'h100000);
  assign T7576 = $signed(31'h2981428b) * $signed(16'h1);
  assign twiddle4_3_95_real = T7579 + T7577;
  assign T7577 = $signed(T7578) / $signed(22'h100000);
  assign T7578 = $signed(31'h3118cdce) * $signed(16'h0);
  assign T7579 = $signed(T7580) / $signed(22'h100000);
  assign T7580 = $signed(31'h290e0660) * $signed(16'h1);
  assign T7581 = T2943[1'h0:1'h0];
  assign T7582 = T2943[1'h1:1'h1];
  assign T7583 = T2943[2'h2:2'h2];
  assign T7584 = T2943[2'h3:2'h3];
  assign T7585 = T2943[3'h4:3'h4];
  assign T7586 = T7803 ? T7681 : T7587;
  assign T7587 = T7680 ? T7634 : T7588;
  assign T7588 = T7633 ? T7611 : T7589;
  assign T7589 = T7610 ? T7600 : T7590;
  assign T7590 = T7599 ? twiddle4_3_97_real : twiddle4_3_96_real;
  assign twiddle4_3_96_real = T7593 + T7591;
  assign T7591 = $signed(T7592) / $signed(22'h100000);
  assign T7592 = $signed(31'h317900d6) * $signed(16'h0);
  assign T7593 = $signed(T7594) / $signed(22'h100000);
  assign T7594 = $signed(31'h2899e64a) * $signed(16'h1);
  assign twiddle4_3_97_real = T7597 + T7595;
  assign T7595 = $signed(T7596) / $signed(22'h100000);
  assign T7596 = $signed(31'h31d82136) * $signed(16'h0);
  assign T7597 = $signed(T7598) / $signed(22'h100000);
  assign T7598 = $signed(31'h2824e4cc) * $signed(16'h1);
  assign T7599 = T2943[1'h0:1'h0];
  assign T7600 = T7609 ? twiddle4_3_99_real : twiddle4_3_98_real;
  assign twiddle4_3_98_real = T7603 + T7601;
  assign T7601 = $signed(T7602) / $signed(22'h100000);
  assign T7602 = $signed(31'h32362cdf) * $signed(16'h0);
  assign T7603 = $signed(T7604) / $signed(22'h100000);
  assign T7604 = $signed(31'h27af0471) * $signed(16'h1);
  assign twiddle4_3_99_real = T7607 + T7605;
  assign T7605 = $signed(T7606) / $signed(22'h100000);
  assign T7606 = $signed(31'h329321c7) * $signed(16'h0);
  assign T7607 = $signed(T7608) / $signed(22'h100000);
  assign T7608 = $signed(31'h273847c7) * $signed(16'h1);
  assign T7609 = T2943[1'h0:1'h0];
  assign T7610 = T2943[1'h1:1'h1];
  assign T7611 = T7632 ? T7622 : T7612;
  assign T7612 = T7621 ? twiddle4_3_101_real : twiddle4_3_100_real;
  assign twiddle4_3_100_real = T7615 + T7613;
  assign T7613 = $signed(T7614) / $signed(22'h100000);
  assign T7614 = $signed(31'h32eefde9) * $signed(16'h0);
  assign T7615 = $signed(T7616) / $signed(22'h100000);
  assign T7616 = $signed(31'h26c0b162) * $signed(16'h1);
  assign twiddle4_3_101_real = T7619 + T7617;
  assign T7617 = $signed(T7618) / $signed(22'h100000);
  assign T7618 = $signed(31'h3349bf48) * $signed(16'h0);
  assign T7619 = $signed(T7620) / $signed(22'h100000);
  assign T7620 = $signed(31'h264843d8) * $signed(16'h1);
  assign T7621 = T2943[1'h0:1'h0];
  assign T7622 = T7631 ? twiddle4_3_103_real : twiddle4_3_102_real;
  assign twiddle4_3_102_real = T7625 + T7623;
  assign T7623 = $signed(T7624) / $signed(22'h100000);
  assign T7624 = $signed(31'h33a363eb) * $signed(16'h0);
  assign T7625 = $signed(T7626) / $signed(22'h100000);
  assign T7626 = $signed(31'h25cf01c7) * $signed(16'h1);
  assign twiddle4_3_103_real = T7629 + T7627;
  assign T7627 = $signed(T7628) / $signed(22'h100000);
  assign T7628 = $signed(31'h33fbe9e2) * $signed(16'h0);
  assign T7629 = $signed(T7630) / $signed(22'h100000);
  assign T7630 = $signed(31'h2554edd0) * $signed(16'h1);
  assign T7631 = T2943[1'h0:1'h0];
  assign T7632 = T2943[1'h1:1'h1];
  assign T7633 = T2943[2'h2:2'h2];
  assign T7634 = T7679 ? T7657 : T7635;
  assign T7635 = T7656 ? T7646 : T7636;
  assign T7636 = T7645 ? twiddle4_3_105_real : twiddle4_3_104_real;
  assign twiddle4_3_104_real = T7639 + T7637;
  assign T7637 = $signed(T7638) / $signed(22'h100000);
  assign T7638 = $signed(31'h34534f40) * $signed(16'h0);
  assign T7639 = $signed(T7640) / $signed(22'h100000);
  assign T7640 = $signed(31'h24da0a99) * $signed(16'h1);
  assign twiddle4_3_105_real = T7643 + T7641;
  assign T7641 = $signed(T7642) / $signed(22'h100000);
  assign T7642 = $signed(31'h34a99221) * $signed(16'h0);
  assign T7643 = $signed(T7644) / $signed(22'h100000);
  assign T7644 = $signed(31'h245e5acc) * $signed(16'h1);
  assign T7645 = T2943[1'h0:1'h0];
  assign T7646 = T7655 ? twiddle4_3_107_real : twiddle4_3_106_real;
  assign twiddle4_3_106_real = T7649 + T7647;
  assign T7647 = $signed(T7648) / $signed(22'h100000);
  assign T7648 = $signed(31'h34feb0a5) * $signed(16'h0);
  assign T7649 = $signed(T7650) / $signed(22'h100000);
  assign T7650 = $signed(31'h23e1e117) * $signed(16'h1);
  assign twiddle4_3_107_real = T7653 + T7651;
  assign T7651 = $signed(T7652) / $signed(22'h100000);
  assign T7652 = $signed(31'h3552a8f4) * $signed(16'h0);
  assign T7653 = $signed(T7654) / $signed(22'h100000);
  assign T7654 = $signed(31'h2364a02e) * $signed(16'h1);
  assign T7655 = T2943[1'h0:1'h0];
  assign T7656 = T2943[1'h1:1'h1];
  assign T7657 = T7678 ? T7668 : T7658;
  assign T7658 = T7667 ? twiddle4_3_109_real : twiddle4_3_108_real;
  assign twiddle4_3_108_real = T7661 + T7659;
  assign T7659 = $signed(T7660) / $signed(22'h100000);
  assign T7660 = $signed(31'h35a5793c) * $signed(16'h0);
  assign T7661 = $signed(T7662) / $signed(22'h100000);
  assign T7662 = $signed(31'h22e69ac7) * $signed(16'h1);
  assign twiddle4_3_109_real = T7665 + T7663;
  assign T7663 = $signed(T7664) / $signed(22'h100000);
  assign T7664 = $signed(31'h35f71fb1) * $signed(16'h0);
  assign T7665 = $signed(T7666) / $signed(22'h100000);
  assign T7666 = $signed(31'h2267d39f) * $signed(16'h1);
  assign T7667 = T2943[1'h0:1'h0];
  assign T7668 = T7677 ? twiddle4_3_111_real : twiddle4_3_110_real;
  assign twiddle4_3_110_real = T7671 + T7669;
  assign T7669 = $signed(T7670) / $signed(22'h100000);
  assign T7670 = $signed(31'h36479a8e) * $signed(16'h0);
  assign T7671 = $signed(T7672) / $signed(22'h100000);
  assign T7672 = $signed(31'h21e84d76) * $signed(16'h1);
  assign twiddle4_3_111_real = T7675 + T7673;
  assign T7673 = $signed(T7674) / $signed(22'h100000);
  assign T7674 = $signed(31'h3696e813) * $signed(16'h0);
  assign T7675 = $signed(T7676) / $signed(22'h100000);
  assign T7676 = $signed(31'h21680b0f) * $signed(16'h1);
  assign T7677 = T2943[1'h0:1'h0];
  assign T7678 = T2943[1'h1:1'h1];
  assign T7679 = T2943[2'h2:2'h2];
  assign T7680 = T2943[2'h3:2'h3];
  assign T7681 = T7802 ? T7740 : T7682;
  assign T7682 = T7739 ? T7709 : T7683;
  assign T7683 = T7708 ? T7694 : T7684;
  assign T7684 = T7693 ? twiddle4_3_113_real : twiddle4_3_112_real;
  assign twiddle4_3_112_real = T7687 + T7685;
  assign T7685 = $signed(T7686) / $signed(22'h100000);
  assign T7686 = $signed(31'h36e5068a) * $signed(16'h0);
  assign T7687 = $signed(T7688) / $signed(22'h100000);
  assign T7688 = $signed(31'h20e70f32) * $signed(16'h1);
  assign twiddle4_3_113_real = T7691 + T7689;
  assign T7689 = $signed(T7690) / $signed(22'h100000);
  assign T7690 = $signed(31'h3731f43f) * $signed(16'h0);
  assign T7691 = $signed(T7692) / $signed(22'h100000);
  assign T7692 = $signed(31'h20655cab) * $signed(16'h1);
  assign T7693 = T2943[1'h0:1'h0];
  assign T7694 = T7707 ? twiddle4_3_115_real : twiddle4_3_114_real;
  assign twiddle4_3_114_real = T7697 + T7695;
  assign T7695 = $signed(T7696) / $signed(22'h100000);
  assign T7696 = $signed(31'h377daf89) * $signed(16'h0);
  assign T7697 = {T7700, T7698};
  assign T7698 = $signed(T7699) / $signed(22'h100000);
  assign T7699 = $signed(30'h1fe2f64b) * $signed(16'h1);
  assign T7700 = T7698[6'h2d:6'h2d];
  assign twiddle4_3_115_real = T7703 + T7701;
  assign T7701 = $signed(T7702) / $signed(22'h100000);
  assign T7702 = $signed(31'h37c836c2) * $signed(16'h0);
  assign T7703 = {T7706, T7704};
  assign T7704 = $signed(T7705) / $signed(22'h100000);
  assign T7705 = $signed(30'h1f5fdee6) * $signed(16'h1);
  assign T7706 = T7704[6'h2d:6'h2d];
  assign T7707 = T2943[1'h0:1'h0];
  assign T7708 = T2943[1'h1:1'h1];
  assign T7709 = T7738 ? T7724 : T7710;
  assign T7710 = T7723 ? twiddle4_3_117_real : twiddle4_3_116_real;
  assign twiddle4_3_116_real = T7713 + T7711;
  assign T7711 = $signed(T7712) / $signed(22'h100000);
  assign T7712 = $signed(31'h3811884c) * $signed(16'h0);
  assign T7713 = {T7716, T7714};
  assign T7714 = $signed(T7715) / $signed(22'h100000);
  assign T7715 = $signed(30'h1edc1952) * $signed(16'h1);
  assign T7716 = T7714[6'h2d:6'h2d];
  assign twiddle4_3_117_real = T7719 + T7717;
  assign T7717 = $signed(T7718) / $signed(22'h100000);
  assign T7718 = $signed(31'h3859a292) * $signed(16'h0);
  assign T7719 = {T7722, T7720};
  assign T7720 = $signed(T7721) / $signed(22'h100000);
  assign T7721 = $signed(30'h1e57a86d) * $signed(16'h1);
  assign T7722 = T7720[6'h2d:6'h2d];
  assign T7723 = T2943[1'h0:1'h0];
  assign T7724 = T7737 ? twiddle4_3_119_real : twiddle4_3_118_real;
  assign twiddle4_3_118_real = T7727 + T7725;
  assign T7725 = $signed(T7726) / $signed(22'h100000);
  assign T7726 = $signed(31'h38a08402) * $signed(16'h0);
  assign T7727 = {T7730, T7728};
  assign T7728 = $signed(T7729) / $signed(22'h100000);
  assign T7729 = $signed(30'h1dd28f14) * $signed(16'h1);
  assign T7730 = T7728[6'h2d:6'h2d];
  assign twiddle4_3_119_real = T7733 + T7731;
  assign T7731 = $signed(T7732) / $signed(22'h100000);
  assign T7732 = $signed(31'h38e62b13) * $signed(16'h0);
  assign T7733 = {T7736, T7734};
  assign T7734 = $signed(T7735) / $signed(22'h100000);
  assign T7735 = $signed(30'h1d4cd02b) * $signed(16'h1);
  assign T7736 = T7734[6'h2d:6'h2d];
  assign T7737 = T2943[1'h0:1'h0];
  assign T7738 = T2943[1'h1:1'h1];
  assign T7739 = T2943[2'h2:2'h2];
  assign T7740 = T7801 ? T7771 : T7741;
  assign T7741 = T7770 ? T7756 : T7742;
  assign T7742 = T7755 ? twiddle4_3_121_real : twiddle4_3_120_real;
  assign twiddle4_3_120_real = T7745 + T7743;
  assign T7743 = $signed(T7744) / $signed(22'h100000);
  assign T7744 = $signed(31'h392a9642) * $signed(16'h0);
  assign T7745 = {T7748, T7746};
  assign T7746 = $signed(T7747) / $signed(22'h100000);
  assign T7747 = $signed(30'h1cc66e99) * $signed(16'h1);
  assign T7748 = T7746[6'h2d:6'h2d];
  assign twiddle4_3_121_real = T7751 + T7749;
  assign T7749 = $signed(T7750) / $signed(22'h100000);
  assign T7750 = $signed(31'h396dc414) * $signed(16'h0);
  assign T7751 = {T7754, T7752};
  assign T7752 = $signed(T7753) / $signed(22'h100000);
  assign T7753 = $signed(30'h1c3f6d47) * $signed(16'h1);
  assign T7754 = T7752[6'h2d:6'h2d];
  assign T7755 = T2943[1'h0:1'h0];
  assign T7756 = T7769 ? twiddle4_3_123_real : twiddle4_3_122_real;
  assign twiddle4_3_122_real = T7759 + T7757;
  assign T7757 = $signed(T7758) / $signed(22'h100000);
  assign T7758 = $signed(31'h39afb313) * $signed(16'h0);
  assign T7759 = {T7762, T7760};
  assign T7760 = $signed(T7761) / $signed(22'h100000);
  assign T7761 = $signed(30'h1bb7cf23) * $signed(16'h1);
  assign T7762 = T7760[6'h2d:6'h2d];
  assign twiddle4_3_123_real = T7765 + T7763;
  assign T7763 = $signed(T7764) / $signed(22'h100000);
  assign T7764 = $signed(31'h39f061d1) * $signed(16'h0);
  assign T7765 = {T7768, T7766};
  assign T7766 = $signed(T7767) / $signed(22'h100000);
  assign T7767 = $signed(30'h1b2f971d) * $signed(16'h1);
  assign T7768 = T7766[6'h2d:6'h2d];
  assign T7769 = T2943[1'h0:1'h0];
  assign T7770 = T2943[1'h1:1'h1];
  assign T7771 = T7800 ? T7786 : T7772;
  assign T7772 = T7785 ? twiddle4_3_125_real : twiddle4_3_124_real;
  assign twiddle4_3_124_real = T7775 + T7773;
  assign T7773 = $signed(T7774) / $signed(22'h100000);
  assign T7774 = $signed(31'h3a2fcee8) * $signed(16'h0);
  assign T7775 = {T7778, T7776};
  assign T7776 = $signed(T7777) / $signed(22'h100000);
  assign T7777 = $signed(30'h1aa6c82b) * $signed(16'h1);
  assign T7778 = T7776[6'h2d:6'h2d];
  assign twiddle4_3_125_real = T7781 + T7779;
  assign T7779 = $signed(T7780) / $signed(22'h100000);
  assign T7780 = $signed(31'h3a6df8f7) * $signed(16'h0);
  assign T7781 = {T7784, T7782};
  assign T7782 = $signed(T7783) / $signed(22'h100000);
  assign T7783 = $signed(30'h1a1d6543) * $signed(16'h1);
  assign T7784 = T7782[6'h2d:6'h2d];
  assign T7785 = T2943[1'h0:1'h0];
  assign T7786 = T7799 ? twiddle4_3_127_real : twiddle4_3_126_real;
  assign twiddle4_3_126_real = T7789 + T7787;
  assign T7787 = $signed(T7788) / $signed(22'h100000);
  assign T7788 = $signed(31'h3aaadea5) * $signed(16'h0);
  assign T7789 = {T7792, T7790};
  assign T7790 = $signed(T7791) / $signed(22'h100000);
  assign T7791 = $signed(30'h19937161) * $signed(16'h1);
  assign T7792 = T7790[6'h2d:6'h2d];
  assign twiddle4_3_127_real = T7795 + T7793;
  assign T7793 = $signed(T7794) / $signed(22'h100000);
  assign T7794 = $signed(31'h3ae67ea1) * $signed(16'h0);
  assign T7795 = {T7798, T7796};
  assign T7796 = $signed(T7797) / $signed(22'h100000);
  assign T7797 = $signed(30'h1908ef81) * $signed(16'h1);
  assign T7798 = T7796[6'h2d:6'h2d];
  assign T7799 = T2943[1'h0:1'h0];
  assign T7800 = T2943[1'h1:1'h1];
  assign T7801 = T2943[2'h2:2'h2];
  assign T7802 = T2943[2'h3:2'h3];
  assign T7803 = T2943[3'h4:3'h4];
  assign T7804 = T2943[3'h5:3'h5];
  assign T7805 = T7395[6'h2e:6'h2e];
  assign T7806 = T2943[3'h6:3'h6];
  assign T7807 = {T8829, T7808};
  assign T7808 = T8828 ? T8367 : T7809;
  assign T7809 = T8366 ? T8080 : T7810;
  assign T7810 = T8079 ? T7937 : T7811;
  assign T7811 = T7936 ? T7874 : T7812;
  assign T7812 = T7873 ? T7843 : T7813;
  assign T7813 = T7842 ? T7828 : T7814;
  assign T7814 = T7827 ? twiddle4_3_129_real : twiddle4_3_128_real;
  assign twiddle4_3_128_real = T7817 + T7815;
  assign T7815 = $signed(T7816) / $signed(22'h100000);
  assign T7816 = $signed(31'h3b20d79e) * $signed(16'h0);
  assign T7817 = {T7820, T7818};
  assign T7818 = $signed(T7819) / $signed(22'h100000);
  assign T7819 = $signed(30'h187de2a6) * $signed(16'h1);
  assign T7820 = T7818[6'h2d:6'h2d];
  assign twiddle4_3_129_real = T7823 + T7821;
  assign T7821 = $signed(T7822) / $signed(22'h100000);
  assign T7822 = $signed(31'h3b59e859) * $signed(16'h0);
  assign T7823 = {T7826, T7824};
  assign T7824 = $signed(T7825) / $signed(22'h100000);
  assign T7825 = $signed(30'h17f24dd3) * $signed(16'h1);
  assign T7826 = T7824[6'h2d:6'h2d];
  assign T7827 = T2943[1'h0:1'h0];
  assign T7828 = T7841 ? twiddle4_3_131_real : twiddle4_3_130_real;
  assign twiddle4_3_130_real = T7831 + T7829;
  assign T7829 = $signed(T7830) / $signed(22'h100000);
  assign T7830 = $signed(31'h3b91af96) * $signed(16'h0);
  assign T7831 = {T7834, T7832};
  assign T7832 = $signed(T7833) / $signed(22'h100000);
  assign T7833 = $signed(30'h1766340f) * $signed(16'h1);
  assign T7834 = T7832[6'h2d:6'h2d];
  assign twiddle4_3_131_real = T7837 + T7835;
  assign T7835 = $signed(T7836) / $signed(22'h100000);
  assign T7836 = $signed(31'h3bc82c1e) * $signed(16'h0);
  assign T7837 = {T7840, T7838};
  assign T7838 = $signed(T7839) / $signed(22'h100000);
  assign T7839 = $signed(30'h16d99863) * $signed(16'h1);
  assign T7840 = T7838[6'h2d:6'h2d];
  assign T7841 = T2943[1'h0:1'h0];
  assign T7842 = T2943[1'h1:1'h1];
  assign T7843 = T7872 ? T7858 : T7844;
  assign T7844 = T7857 ? twiddle4_3_133_real : twiddle4_3_132_real;
  assign twiddle4_3_132_real = T7847 + T7845;
  assign T7845 = $signed(T7846) / $signed(22'h100000);
  assign T7846 = $signed(31'h3bfd5cc4) * $signed(16'h0);
  assign T7847 = {T7850, T7848};
  assign T7848 = $signed(T7849) / $signed(22'h100000);
  assign T7849 = $signed(30'h164c7ddd) * $signed(16'h1);
  assign T7850 = T7848[6'h2d:6'h2d];
  assign twiddle4_3_133_real = T7853 + T7851;
  assign T7851 = $signed(T7852) / $signed(22'h100000);
  assign T7852 = $signed(31'h3c31405f) * $signed(16'h0);
  assign T7853 = {T7856, T7854};
  assign T7854 = $signed(T7855) / $signed(22'h100000);
  assign T7855 = $signed(30'h15bee78b) * $signed(16'h1);
  assign T7856 = T7854[6'h2d:6'h2d];
  assign T7857 = T2943[1'h0:1'h0];
  assign T7858 = T7871 ? twiddle4_3_135_real : twiddle4_3_134_real;
  assign twiddle4_3_134_real = T7861 + T7859;
  assign T7859 = $signed(T7860) / $signed(22'h100000);
  assign T7860 = $signed(31'h3c63d5d0) * $signed(16'h0);
  assign T7861 = {T7864, T7862};
  assign T7862 = $signed(T7863) / $signed(22'h100000);
  assign T7863 = $signed(30'h1530d880) * $signed(16'h1);
  assign T7864 = T7862[6'h2d:6'h2d];
  assign twiddle4_3_135_real = T7867 + T7865;
  assign T7865 = $signed(T7866) / $signed(22'h100000);
  assign T7866 = $signed(31'h3c951bff) * $signed(16'h0);
  assign T7867 = {T7870, T7868};
  assign T7868 = $signed(T7869) / $signed(22'h100000);
  assign T7869 = $signed(30'h14a253d1) * $signed(16'h1);
  assign T7870 = T7868[6'h2d:6'h2d];
  assign T7871 = T2943[1'h0:1'h0];
  assign T7872 = T2943[1'h1:1'h1];
  assign T7873 = T2943[2'h2:2'h2];
  assign T7874 = T7935 ? T7905 : T7875;
  assign T7875 = T7904 ? T7890 : T7876;
  assign T7876 = T7889 ? twiddle4_3_137_real : twiddle4_3_136_real;
  assign twiddle4_3_136_real = T7879 + T7877;
  assign T7877 = $signed(T7878) / $signed(22'h100000);
  assign T7878 = $signed(31'h3cc511d8) * $signed(16'h0);
  assign T7879 = {T7882, T7880};
  assign T7880 = $signed(T7881) / $signed(22'h100000);
  assign T7881 = $signed(30'h14135c94) * $signed(16'h1);
  assign T7882 = T7880[6'h2d:6'h2d];
  assign twiddle4_3_137_real = T7885 + T7883;
  assign T7883 = $signed(T7884) / $signed(22'h100000);
  assign T7884 = $signed(31'h3cf3b653) * $signed(16'h0);
  assign T7885 = {T7888, T7886};
  assign T7886 = $signed(T7887) / $signed(22'h100000);
  assign T7887 = $signed(30'h1383f5e3) * $signed(16'h1);
  assign T7888 = T7886[6'h2d:6'h2d];
  assign T7889 = T2943[1'h0:1'h0];
  assign T7890 = T7903 ? twiddle4_3_139_real : twiddle4_3_138_real;
  assign twiddle4_3_138_real = T7893 + T7891;
  assign T7891 = $signed(T7892) / $signed(22'h100000);
  assign T7892 = $signed(31'h3d21086c) * $signed(16'h0);
  assign T7893 = {T7896, T7894};
  assign T7894 = $signed(T7895) / $signed(22'h100000);
  assign T7895 = $signed(30'h12f422da) * $signed(16'h1);
  assign T7896 = T7894[6'h2d:6'h2d];
  assign twiddle4_3_139_real = T7899 + T7897;
  assign T7897 = $signed(T7898) / $signed(22'h100000);
  assign T7898 = $signed(31'h3d4d0727) * $signed(16'h0);
  assign T7899 = {T7902, T7900};
  assign T7900 = $signed(T7901) / $signed(22'h100000);
  assign T7901 = $signed(30'h1263e699) * $signed(16'h1);
  assign T7902 = T7900[6'h2d:6'h2d];
  assign T7903 = T2943[1'h0:1'h0];
  assign T7904 = T2943[1'h1:1'h1];
  assign T7905 = T7934 ? T7920 : T7906;
  assign T7906 = T7919 ? twiddle4_3_141_real : twiddle4_3_140_real;
  assign twiddle4_3_140_real = T7909 + T7907;
  assign T7907 = $signed(T7908) / $signed(22'h100000);
  assign T7908 = $signed(31'h3d77b191) * $signed(16'h0);
  assign T7909 = {T7912, T7910};
  assign T7910 = $signed(T7911) / $signed(22'h100000);
  assign T7911 = $signed(30'h11d3443f) * $signed(16'h1);
  assign T7912 = T7910[6'h2d:6'h2d];
  assign twiddle4_3_141_real = T7915 + T7913;
  assign T7913 = $signed(T7914) / $signed(22'h100000);
  assign T7914 = $signed(31'h3da106bd) * $signed(16'h0);
  assign T7915 = {T7918, T7916};
  assign T7916 = $signed(T7917) / $signed(22'h100000);
  assign T7917 = $signed(30'h11423eef) * $signed(16'h1);
  assign T7918 = T7916[6'h2d:6'h2d];
  assign T7919 = T2943[1'h0:1'h0];
  assign T7920 = T7933 ? twiddle4_3_143_real : twiddle4_3_142_real;
  assign twiddle4_3_142_real = T7923 + T7921;
  assign T7921 = $signed(T7922) / $signed(22'h100000);
  assign T7922 = $signed(31'h3dc905c4) * $signed(16'h0);
  assign T7923 = {T7926, T7924};
  assign T7924 = $signed(T7925) / $signed(22'h100000);
  assign T7925 = $signed(30'h10b0d9cf) * $signed(16'h1);
  assign T7926 = T7924[6'h2d:6'h2d];
  assign twiddle4_3_143_real = T7929 + T7927;
  assign T7927 = $signed(T7928) / $signed(22'h100000);
  assign T7928 = $signed(31'h3defadca) * $signed(16'h0);
  assign T7929 = {T7932, T7930};
  assign T7930 = $signed(T7931) / $signed(22'h100000);
  assign T7931 = $signed(30'h101f1806) * $signed(16'h1);
  assign T7932 = T7930[6'h2d:6'h2d];
  assign T7933 = T2943[1'h0:1'h0];
  assign T7934 = T2943[1'h1:1'h1];
  assign T7935 = T2943[2'h2:2'h2];
  assign T7936 = T2943[2'h3:2'h3];
  assign T7937 = T8078 ? T8008 : T7938;
  assign T7938 = T8007 ? T7973 : T7939;
  assign T7939 = T7972 ? T7956 : T7940;
  assign T7940 = T7955 ? twiddle4_3_145_real : twiddle4_3_144_real;
  assign twiddle4_3_144_real = T7943 + T7941;
  assign T7941 = $signed(T7942) / $signed(22'h100000);
  assign T7942 = $signed(31'h3e14fdf7) * $signed(16'h0);
  assign T7943 = {T7946, T7944};
  assign T7944 = $signed(T7945) / $signed(22'h100000);
  assign T7945 = $signed(29'hf8cfcbd) * $signed(16'h1);
  assign T7946 = T7947 ? 2'h3 : 2'h0;
  assign T7947 = T7944[6'h2c:6'h2c];
  assign twiddle4_3_145_real = T7950 + T7948;
  assign T7948 = $signed(T7949) / $signed(22'h100000);
  assign T7949 = $signed(31'h3e38f57c) * $signed(16'h0);
  assign T7950 = {T7953, T7951};
  assign T7951 = $signed(T7952) / $signed(22'h100000);
  assign T7952 = $signed(29'hefa8b1f) * $signed(16'h1);
  assign T7953 = T7954 ? 2'h3 : 2'h0;
  assign T7954 = T7951[6'h2c:6'h2c];
  assign T7955 = T2943[1'h0:1'h0];
  assign T7956 = T7971 ? twiddle4_3_147_real : twiddle4_3_146_real;
  assign twiddle4_3_146_real = T7959 + T7957;
  assign T7957 = $signed(T7958) / $signed(22'h100000);
  assign T7958 = $signed(31'h3e5b9392) * $signed(16'h0);
  assign T7959 = {T7962, T7960};
  assign T7960 = $signed(T7961) / $signed(22'h100000);
  assign T7961 = $signed(29'he67c659) * $signed(16'h1);
  assign T7962 = T7963 ? 2'h3 : 2'h0;
  assign T7963 = T7960[6'h2c:6'h2c];
  assign twiddle4_3_147_real = T7966 + T7964;
  assign T7964 = $signed(T7965) / $signed(22'h100000);
  assign T7965 = $signed(31'h3e7cd778) * $signed(16'h0);
  assign T7966 = {T7969, T7967};
  assign T7967 = $signed(T7968) / $signed(22'h100000);
  assign T7968 = $signed(29'hdd4b19a) * $signed(16'h1);
  assign T7969 = T7970 ? 2'h3 : 2'h0;
  assign T7970 = T7967[6'h2c:6'h2c];
  assign T7971 = T2943[1'h0:1'h0];
  assign T7972 = T2943[1'h1:1'h1];
  assign T7973 = T8006 ? T7990 : T7974;
  assign T7974 = T7989 ? twiddle4_3_149_real : twiddle4_3_148_real;
  assign twiddle4_3_148_real = T7977 + T7975;
  assign T7975 = $signed(T7976) / $signed(22'h100000);
  assign T7976 = $signed(31'h3e9cc076) * $signed(16'h0);
  assign T7977 = {T7980, T7978};
  assign T7978 = $signed(T7979) / $signed(22'h100000);
  assign T7979 = $signed(29'hd415012) * $signed(16'h1);
  assign T7980 = T7981 ? 2'h3 : 2'h0;
  assign T7981 = T7978[6'h2c:6'h2c];
  assign twiddle4_3_149_real = T7984 + T7982;
  assign T7982 = $signed(T7983) / $signed(22'h100000);
  assign T7983 = $signed(31'h3ebb4dda) * $signed(16'h0);
  assign T7984 = {T7987, T7985};
  assign T7985 = $signed(T7986) / $signed(22'h100000);
  assign T7986 = $signed(29'hcada4f4) * $signed(16'h1);
  assign T7987 = T7988 ? 2'h3 : 2'h0;
  assign T7988 = T7985[6'h2c:6'h2c];
  assign T7989 = T2943[1'h0:1'h0];
  assign T7990 = T8005 ? twiddle4_3_151_real : twiddle4_3_150_real;
  assign twiddle4_3_150_real = T7993 + T7991;
  assign T7991 = $signed(T7992) / $signed(22'h100000);
  assign T7992 = $signed(31'h3ed87efb) * $signed(16'h0);
  assign T7993 = {T7996, T7994};
  assign T7994 = $signed(T7995) / $signed(22'h100000);
  assign T7995 = $signed(29'hc19b374) * $signed(16'h1);
  assign T7996 = T7997 ? 2'h3 : 2'h0;
  assign T7997 = T7994[6'h2c:6'h2c];
  assign twiddle4_3_151_real = T8000 + T7998;
  assign T7998 = $signed(T7999) / $signed(22'h100000);
  assign T7999 = $signed(31'h3ef45338) * $signed(16'h0);
  assign T8000 = {T8003, T8001};
  assign T8001 = $signed(T8002) / $signed(22'h100000);
  assign T8002 = $signed(29'hb857ec6) * $signed(16'h1);
  assign T8003 = T8004 ? 2'h3 : 2'h0;
  assign T8004 = T8001[6'h2c:6'h2c];
  assign T8005 = T2943[1'h0:1'h0];
  assign T8006 = T2943[1'h1:1'h1];
  assign T8007 = T2943[2'h2:2'h2];
  assign T8008 = T8077 ? T8043 : T8009;
  assign T8009 = T8042 ? T8026 : T8010;
  assign T8010 = T8025 ? twiddle4_3_153_real : twiddle4_3_152_real;
  assign twiddle4_3_152_real = T8013 + T8011;
  assign T8011 = $signed(T8012) / $signed(22'h100000);
  assign T8012 = $signed(31'h3f0ec9f4) * $signed(16'h0);
  assign T8013 = {T8016, T8014};
  assign T8014 = $signed(T8015) / $signed(22'h100000);
  assign T8015 = $signed(29'haf10a22) * $signed(16'h1);
  assign T8016 = T8017 ? 2'h3 : 2'h0;
  assign T8017 = T8014[6'h2c:6'h2c];
  assign twiddle4_3_153_real = T8020 + T8018;
  assign T8018 = $signed(T8019) / $signed(22'h100000);
  assign T8019 = $signed(31'h3f27e29f) * $signed(16'h0);
  assign T8020 = {T8023, T8021};
  assign T8021 = $signed(T8022) / $signed(22'h100000);
  assign T8022 = $signed(29'ha5c58bf) * $signed(16'h1);
  assign T8023 = T8024 ? 2'h3 : 2'h0;
  assign T8024 = T8021[6'h2c:6'h2c];
  assign T8025 = T2943[1'h0:1'h0];
  assign T8026 = T8041 ? twiddle4_3_155_real : twiddle4_3_154_real;
  assign twiddle4_3_154_real = T8029 + T8027;
  assign T8027 = $signed(T8028) / $signed(22'h100000);
  assign T8028 = $signed(31'h3f3f9cab) * $signed(16'h0);
  assign T8029 = {T8032, T8030};
  assign T8030 = $signed(T8031) / $signed(22'h100000);
  assign T8031 = $signed(29'h9c76dd8) * $signed(16'h1);
  assign T8032 = T8033 ? 2'h3 : 2'h0;
  assign T8033 = T8030[6'h2c:6'h2c];
  assign twiddle4_3_155_real = T8036 + T8034;
  assign T8034 = $signed(T8035) / $signed(22'h100000);
  assign T8035 = $signed(31'h3f55f796) * $signed(16'h0);
  assign T8036 = {T8039, T8037};
  assign T8037 = $signed(T8038) / $signed(22'h100000);
  assign T8038 = $signed(29'h9324ca6) * $signed(16'h1);
  assign T8039 = T8040 ? 2'h3 : 2'h0;
  assign T8040 = T8037[6'h2c:6'h2c];
  assign T8041 = T2943[1'h0:1'h0];
  assign T8042 = T2943[1'h1:1'h1];
  assign T8043 = T8076 ? T8060 : T8044;
  assign T8044 = T8059 ? twiddle4_3_157_real : twiddle4_3_156_real;
  assign twiddle4_3_156_real = T8047 + T8045;
  assign T8045 = $signed(T8046) / $signed(22'h100000);
  assign T8046 = $signed(31'h3f6af2e3) * $signed(16'h0);
  assign T8047 = {T8050, T8048};
  assign T8048 = $signed(T8049) / $signed(22'h100000);
  assign T8049 = $signed(29'h89cf867) * $signed(16'h1);
  assign T8050 = T8051 ? 2'h3 : 2'h0;
  assign T8051 = T8048[6'h2c:6'h2c];
  assign twiddle4_3_157_real = T8054 + T8052;
  assign T8052 = $signed(T8053) / $signed(22'h100000);
  assign T8053 = $signed(31'h3f7e8e1e) * $signed(16'h0);
  assign T8054 = {T8057, T8055};
  assign T8055 = $signed(T8056) / $signed(22'h100000);
  assign T8056 = $signed(29'h8077456) * $signed(16'h1);
  assign T8057 = T8058 ? 2'h3 : 2'h0;
  assign T8058 = T8055[6'h2c:6'h2c];
  assign T8059 = T2943[1'h0:1'h0];
  assign T8060 = T8075 ? twiddle4_3_159_real : twiddle4_3_158_real;
  assign twiddle4_3_158_real = T8063 + T8061;
  assign T8061 = $signed(T8062) / $signed(22'h100000);
  assign T8062 = $signed(31'h3f90c8d9) * $signed(16'h0);
  assign T8063 = {T8066, T8064};
  assign T8064 = $signed(T8065) / $signed(22'h100000);
  assign T8065 = $signed(28'h771c3b2) * $signed(16'h1);
  assign T8066 = T8067 ? 3'h7 : 3'h0;
  assign T8067 = T8064[6'h2b:6'h2b];
  assign twiddle4_3_159_real = T8070 + T8068;
  assign T8068 = $signed(T8069) / $signed(22'h100000);
  assign T8069 = $signed(31'h3fa1a2b1) * $signed(16'h0);
  assign T8070 = {T8073, T8071};
  assign T8071 = $signed(T8072) / $signed(22'h100000);
  assign T8072 = $signed(28'h6dbe9bb) * $signed(16'h1);
  assign T8073 = T8074 ? 3'h7 : 3'h0;
  assign T8074 = T8071[6'h2b:6'h2b];
  assign T8075 = T2943[1'h0:1'h0];
  assign T8076 = T2943[1'h1:1'h1];
  assign T8077 = T2943[2'h2:2'h2];
  assign T8078 = T2943[2'h3:2'h3];
  assign T8079 = T2943[3'h4:3'h4];
  assign T8080 = T8365 ? T8223 : T8081;
  assign T8081 = T8222 ? T8152 : T8082;
  assign T8082 = T8151 ? T8117 : T8083;
  assign T8083 = T8116 ? T8100 : T8084;
  assign T8084 = T8099 ? twiddle4_3_161_real : twiddle4_3_160_real;
  assign twiddle4_3_160_real = T8087 + T8085;
  assign T8085 = $signed(T8086) / $signed(22'h100000);
  assign T8086 = $signed(31'h3fb11b47) * $signed(16'h0);
  assign T8087 = {T8090, T8088};
  assign T8088 = $signed(T8089) / $signed(22'h100000);
  assign T8089 = $signed(28'h645e9af) * $signed(16'h1);
  assign T8090 = T8091 ? 3'h7 : 3'h0;
  assign T8091 = T8088[6'h2b:6'h2b];
  assign twiddle4_3_161_real = T8094 + T8092;
  assign T8092 = $signed(T8093) / $signed(22'h100000);
  assign T8093 = $signed(31'h3fbf3245) * $signed(16'h0);
  assign T8094 = {T8097, T8095};
  assign T8095 = $signed(T8096) / $signed(22'h100000);
  assign T8096 = $signed(28'h5afc6cf) * $signed(16'h1);
  assign T8097 = T8098 ? 3'h7 : 3'h0;
  assign T8098 = T8095[6'h2b:6'h2b];
  assign T8099 = T2943[1'h0:1'h0];
  assign T8100 = T8115 ? twiddle4_3_163_real : twiddle4_3_162_real;
  assign twiddle4_3_162_real = T8103 + T8101;
  assign T8101 = $signed(T8102) / $signed(22'h100000);
  assign T8102 = $signed(31'h3fcbe75e) * $signed(16'h0);
  assign T8103 = {T8106, T8104};
  assign T8104 = $signed(T8105) / $signed(22'h100000);
  assign T8105 = $signed(28'h519845e) * $signed(16'h1);
  assign T8106 = T8107 ? 3'h7 : 3'h0;
  assign T8107 = T8104[6'h2b:6'h2b];
  assign twiddle4_3_163_real = T8110 + T8108;
  assign T8108 = $signed(T8109) / $signed(22'h100000);
  assign T8109 = $signed(31'h3fd73a4a) * $signed(16'h0);
  assign T8110 = {T8113, T8111};
  assign T8111 = $signed(T8112) / $signed(22'h100000);
  assign T8112 = $signed(28'h483259d) * $signed(16'h1);
  assign T8113 = T8114 ? 3'h7 : 3'h0;
  assign T8114 = T8111[6'h2b:6'h2b];
  assign T8115 = T2943[1'h0:1'h0];
  assign T8116 = T2943[1'h1:1'h1];
  assign T8117 = T8150 ? T8134 : T8118;
  assign T8118 = T8133 ? twiddle4_3_165_real : twiddle4_3_164_real;
  assign twiddle4_3_164_real = T8121 + T8119;
  assign T8119 = $signed(T8120) / $signed(22'h100000);
  assign T8120 = $signed(31'h3fe12acb) * $signed(16'h0);
  assign T8121 = {T8124, T8122};
  assign T8122 = $signed(T8123) / $signed(22'h100000);
  assign T8123 = $signed(27'h3ecadcf) * $signed(16'h1);
  assign T8124 = T8125 ? 4'hf : 4'h0;
  assign T8125 = T8122[6'h2a:6'h2a];
  assign twiddle4_3_165_real = T8128 + T8126;
  assign T8126 = $signed(T8127) / $signed(22'h100000);
  assign T8127 = $signed(31'h3fe9b8a9) * $signed(16'h0);
  assign T8128 = {T8131, T8129};
  assign T8129 = $signed(T8130) / $signed(22'h100000);
  assign T8130 = $signed(27'h3562037) * $signed(16'h1);
  assign T8131 = T8132 ? 4'hf : 4'h0;
  assign T8132 = T8129[6'h2a:6'h2a];
  assign T8133 = T2943[1'h0:1'h0];
  assign T8134 = T8149 ? twiddle4_3_167_real : twiddle4_3_166_real;
  assign twiddle4_3_166_real = T8137 + T8135;
  assign T8135 = $signed(T8136) / $signed(22'h100000);
  assign T8136 = $signed(31'h3ff0e3b5) * $signed(16'h0);
  assign T8137 = {T8140, T8138};
  assign T8138 = $signed(T8139) / $signed(22'h100000);
  assign T8139 = $signed(27'h2bf801a) * $signed(16'h1);
  assign T8140 = T8141 ? 4'hf : 4'h0;
  assign T8141 = T8138[6'h2a:6'h2a];
  assign twiddle4_3_167_real = T8144 + T8142;
  assign T8142 = $signed(T8143) / $signed(22'h100000);
  assign T8143 = $signed(31'h3ff6abc8) * $signed(16'h0);
  assign T8144 = {T8147, T8145};
  assign T8145 = $signed(T8146) / $signed(22'h100000);
  assign T8146 = $signed(27'h228d0bb) * $signed(16'h1);
  assign T8147 = T8148 ? 4'hf : 4'h0;
  assign T8148 = T8145[6'h2a:6'h2a];
  assign T8149 = T2943[1'h0:1'h0];
  assign T8150 = T2943[1'h1:1'h1];
  assign T8151 = T2943[2'h2:2'h2];
  assign T8152 = T8221 ? T8187 : T8153;
  assign T8153 = T8186 ? T8170 : T8154;
  assign T8154 = T8169 ? twiddle4_3_169_real : twiddle4_3_168_real;
  assign twiddle4_3_168_real = T8157 + T8155;
  assign T8155 = $signed(T8156) / $signed(22'h100000);
  assign T8156 = $signed(31'h3ffb10c1) * $signed(16'h0);
  assign T8157 = {T8160, T8158};
  assign T8158 = $signed(T8159) / $signed(22'h100000);
  assign T8159 = $signed(26'h192155f) * $signed(16'h1);
  assign T8160 = T8161 ? 5'h1f : 5'h0;
  assign T8161 = T8158[6'h29:6'h29];
  assign twiddle4_3_169_real = T8164 + T8162;
  assign T8162 = $signed(T8163) / $signed(22'h100000);
  assign T8163 = $signed(31'h3ffe1287) * $signed(16'h0);
  assign T8164 = {T8167, T8165};
  assign T8165 = $signed(T8166) / $signed(22'h100000);
  assign T8166 = $signed(25'hfb514b) * $signed(16'h1);
  assign T8167 = T8168 ? 6'h3f : 6'h0;
  assign T8168 = T8165[6'h28:6'h28];
  assign T8169 = T2943[1'h0:1'h0];
  assign T8170 = T8185 ? twiddle4_3_171_real : twiddle4_3_170_real;
  assign twiddle4_3_170_real = T8173 + T8171;
  assign T8171 = $signed(T8172) / $signed(22'h100000);
  assign T8172 = $signed(31'h3fffb10b) * $signed(16'h0);
  assign T8173 = {T8176, T8174};
  assign T8174 = $signed(T8175) / $signed(22'h100000);
  assign T8175 = $signed(24'h6487c3) * $signed(16'h1);
  assign T8176 = T8177 ? 7'h7f : 7'h0;
  assign T8177 = T8174[6'h27:6'h27];
  assign twiddle4_3_171_real = T8180 + T8178;
  assign T8178 = $signed(T8179) / $signed(22'h100000);
  assign T8179 = $signed(31'h3fffec42) * $signed(16'h0);
  assign T8180 = {T8183, T8181};
  assign T8181 = $signed(T8182) / $signed(22'h100000);
  assign T8182 = $signed(23'h4dbc0f) * $signed(16'h1);
  assign T8183 = T8184 ? 8'hff : 8'h0;
  assign T8184 = T8181[6'h26:6'h26];
  assign T8185 = T2943[1'h0:1'h0];
  assign T8186 = T2943[1'h1:1'h1];
  assign T8187 = T8220 ? T8204 : T8188;
  assign T8188 = T8203 ? twiddle4_3_173_real : twiddle4_3_172_real;
  assign twiddle4_3_172_real = T8191 + T8189;
  assign T8189 = $signed(T8190) / $signed(22'h100000);
  assign T8190 = $signed(31'h3ffec42d) * $signed(16'h0);
  assign T8191 = {T8194, T8192};
  assign T8192 = $signed(T8193) / $signed(22'h100000);
  assign T8193 = $signed(25'h136f171) * $signed(16'h1);
  assign T8194 = T8195 ? 6'h3f : 6'h0;
  assign T8195 = T8192[6'h28:6'h28];
  assign twiddle4_3_173_real = T8198 + T8196;
  assign T8196 = $signed(T8197) / $signed(22'h100000);
  assign T8197 = $signed(31'h3ffc38d0) * $signed(16'h0);
  assign T8198 = {T8201, T8199};
  assign T8199 = $signed(T8200) / $signed(22'h100000);
  assign T8200 = $signed(26'h2a02b2e) * $signed(16'h1);
  assign T8201 = T8202 ? 5'h1f : 5'h0;
  assign T8202 = T8199[6'h29:6'h29];
  assign T8203 = T2943[1'h0:1'h0];
  assign T8204 = T8219 ? twiddle4_3_175_real : twiddle4_3_174_real;
  assign twiddle4_3_174_real = T8207 + T8205;
  assign T8205 = $signed(T8206) / $signed(22'h100000);
  assign T8206 = $signed(31'h3ff84a3b) * $signed(16'h0);
  assign T8207 = {T8210, T8208};
  assign T8208 = $signed(T8209) / $signed(22'h100000);
  assign T8209 = $signed(26'h2096c8d) * $signed(16'h1);
  assign T8210 = T8211 ? 5'h1f : 5'h0;
  assign T8211 = T8208[6'h29:6'h29];
  assign twiddle4_3_175_real = T8214 + T8212;
  assign T8212 = $signed(T8213) / $signed(22'h100000);
  assign T8213 = $signed(31'h3ff2f884) * $signed(16'h0);
  assign T8214 = {T8217, T8215};
  assign T8215 = $signed(T8216) / $signed(22'h100000);
  assign T8216 = $signed(27'h572b8d3) * $signed(16'h1);
  assign T8217 = T8218 ? 4'hf : 4'h0;
  assign T8218 = T8215[6'h2a:6'h2a];
  assign T8219 = T2943[1'h0:1'h0];
  assign T8220 = T2943[1'h1:1'h1];
  assign T8221 = T2943[2'h2:2'h2];
  assign T8222 = T2943[2'h3:2'h3];
  assign T8223 = T8364 ? T8294 : T8224;
  assign T8224 = T8293 ? T8259 : T8225;
  assign T8225 = T8258 ? T8242 : T8226;
  assign T8226 = T8241 ? twiddle4_3_177_real : twiddle4_3_176_real;
  assign twiddle4_3_176_real = T8229 + T8227;
  assign T8227 = $signed(T8228) / $signed(22'h100000);
  assign T8228 = $signed(31'h3fec43c6) * $signed(16'h0);
  assign T8229 = {T8232, T8230};
  assign T8230 = $signed(T8231) / $signed(22'h100000);
  assign T8231 = $signed(27'h4dc1342) * $signed(16'h1);
  assign T8232 = T8233 ? 4'hf : 4'h0;
  assign T8233 = T8230[6'h2a:6'h2a];
  assign twiddle4_3_177_real = T8236 + T8234;
  assign T8234 = $signed(T8235) / $signed(22'h100000);
  assign T8235 = $signed(31'h3fe42c29) * $signed(16'h0);
  assign T8236 = {T8239, T8237};
  assign T8237 = $signed(T8238) / $signed(22'h100000);
  assign T8238 = $signed(27'h4457f21) * $signed(16'h1);
  assign T8239 = T8240 ? 4'hf : 4'h0;
  assign T8240 = T8237[6'h2a:6'h2a];
  assign T8241 = T2943[1'h0:1'h0];
  assign T8242 = T8257 ? twiddle4_3_179_real : twiddle4_3_178_real;
  assign twiddle4_3_178_real = T8245 + T8243;
  assign T8243 = $signed(T8244) / $signed(22'h100000);
  assign T8244 = $signed(31'h3fdab1d9) * $signed(16'h0);
  assign T8245 = {T8248, T8246};
  assign T8246 = $signed(T8247) / $signed(22'h100000);
  assign T8247 = $signed(28'hbaeffb3) * $signed(16'h1);
  assign T8248 = T8249 ? 3'h7 : 3'h0;
  assign T8249 = T8246[6'h2b:6'h2b];
  assign twiddle4_3_179_real = T8252 + T8250;
  assign T8250 = $signed(T8251) / $signed(22'h100000);
  assign T8251 = $signed(31'h3fcfd50a) * $signed(16'h0);
  assign T8252 = {T8255, T8253};
  assign T8253 = $signed(T8254) / $signed(22'h100000);
  assign T8254 = $signed(28'hb18983c) * $signed(16'h1);
  assign T8255 = T8256 ? 3'h7 : 3'h0;
  assign T8256 = T8253[6'h2b:6'h2b];
  assign T8257 = T2943[1'h0:1'h0];
  assign T8258 = T2943[1'h1:1'h1];
  assign T8259 = T8292 ? T8276 : T8260;
  assign T8260 = T8275 ? twiddle4_3_181_real : twiddle4_3_180_real;
  assign twiddle4_3_180_real = T8263 + T8261;
  assign T8261 = $signed(T8262) / $signed(22'h100000);
  assign T8262 = $signed(31'h3fc395f9) * $signed(16'h0);
  assign T8263 = {T8266, T8264};
  assign T8264 = $signed(T8265) / $signed(22'h100000);
  assign T8265 = $signed(28'ha824bfe) * $signed(16'h1);
  assign T8266 = T8267 ? 3'h7 : 3'h0;
  assign T8267 = T8264[6'h2b:6'h2b];
  assign twiddle4_3_181_real = T8270 + T8268;
  assign T8268 = $signed(T8269) / $signed(22'h100000);
  assign T8269 = $signed(31'h3fb5f4ea) * $signed(16'h0);
  assign T8270 = {T8273, T8271};
  assign T8271 = $signed(T8272) / $signed(22'h100000);
  assign T8272 = $signed(28'h9ec1e3c) * $signed(16'h1);
  assign T8273 = T8274 ? 3'h7 : 3'h0;
  assign T8274 = T8271[6'h2b:6'h2b];
  assign T8275 = T2943[1'h0:1'h0];
  assign T8276 = T8291 ? twiddle4_3_183_real : twiddle4_3_182_real;
  assign twiddle4_3_182_real = T8279 + T8277;
  assign T8277 = $signed(T8278) / $signed(22'h100000);
  assign T8278 = $signed(31'h3fa6f228) * $signed(16'h0);
  assign T8279 = {T8282, T8280};
  assign T8280 = $signed(T8281) / $signed(22'h100000);
  assign T8281 = $signed(28'h9561237) * $signed(16'h1);
  assign T8282 = T8283 ? 3'h7 : 3'h0;
  assign T8283 = T8280[6'h2b:6'h2b];
  assign twiddle4_3_183_real = T8286 + T8284;
  assign T8284 = $signed(T8285) / $signed(22'h100000);
  assign T8285 = $signed(31'h3f968e07) * $signed(16'h0);
  assign T8286 = {T8289, T8287};
  assign T8287 = $signed(T8288) / $signed(22'h100000);
  assign T8288 = $signed(28'h8c02b32) * $signed(16'h1);
  assign T8289 = T8290 ? 3'h7 : 3'h0;
  assign T8290 = T8287[6'h2b:6'h2b];
  assign T8291 = T2943[1'h0:1'h0];
  assign T8292 = T2943[1'h1:1'h1];
  assign T8293 = T2943[2'h2:2'h2];
  assign T8294 = T8363 ? T8329 : T8295;
  assign T8295 = T8328 ? T8312 : T8296;
  assign T8296 = T8311 ? twiddle4_3_185_real : twiddle4_3_184_real;
  assign twiddle4_3_184_real = T8299 + T8297;
  assign T8297 = $signed(T8298) / $signed(22'h100000);
  assign T8298 = $signed(31'h3f84c8e1) * $signed(16'h0);
  assign T8299 = {T8302, T8300};
  assign T8300 = $signed(T8301) / $signed(22'h100000);
  assign T8301 = $signed(28'h82a6c6b) * $signed(16'h1);
  assign T8302 = T8303 ? 3'h7 : 3'h0;
  assign T8303 = T8300[6'h2b:6'h2b];
  assign twiddle4_3_185_real = T8306 + T8304;
  assign T8304 = $signed(T8305) / $signed(22'h100000);
  assign T8305 = $signed(31'h3f71a31a) * $signed(16'h0);
  assign T8306 = {T8309, T8307};
  assign T8307 = $signed(T8308) / $signed(22'h100000);
  assign T8308 = $signed(29'h1794d922) * $signed(16'h1);
  assign T8309 = T8310 ? 2'h3 : 2'h0;
  assign T8310 = T8307[6'h2c:6'h2c];
  assign T8311 = T2943[1'h0:1'h0];
  assign T8312 = T8327 ? twiddle4_3_187_real : twiddle4_3_186_real;
  assign twiddle4_3_186_real = T8315 + T8313;
  assign T8313 = $signed(T8314) / $signed(22'h100000);
  assign T8314 = $signed(31'h3f5d1d1c) * $signed(16'h0);
  assign T8315 = {T8318, T8316};
  assign T8316 = $signed(T8317) / $signed(22'h100000);
  assign T8317 = $signed(29'h16ff7496) * $signed(16'h1);
  assign T8318 = T8319 ? 2'h3 : 2'h0;
  assign T8319 = T8316[6'h2c:6'h2c];
  assign twiddle4_3_187_real = T8322 + T8320;
  assign T8320 = $signed(T8321) / $signed(22'h100000);
  assign T8321 = $signed(31'h3f473758) * $signed(16'h0);
  assign T8322 = {T8325, T8323};
  assign T8323 = $signed(T8324) / $signed(22'h100000);
  assign T8324 = $signed(29'h166a4204) * $signed(16'h1);
  assign T8325 = T8326 ? 2'h3 : 2'h0;
  assign T8326 = T8323[6'h2c:6'h2c];
  assign T8327 = T2943[1'h0:1'h0];
  assign T8328 = T2943[1'h1:1'h1];
  assign T8329 = T8362 ? T8346 : T8330;
  assign T8330 = T8345 ? twiddle4_3_189_real : twiddle4_3_188_real;
  assign twiddle4_3_188_real = T8333 + T8331;
  assign T8331 = $signed(T8332) / $signed(22'h100000);
  assign T8332 = $signed(31'h3f2ff249) * $signed(16'h0);
  assign T8333 = {T8336, T8334};
  assign T8334 = $signed(T8335) / $signed(22'h100000);
  assign T8335 = $signed(29'h15d544a8) * $signed(16'h1);
  assign T8336 = T8337 ? 2'h3 : 2'h0;
  assign T8337 = T8334[6'h2c:6'h2c];
  assign twiddle4_3_189_real = T8340 + T8338;
  assign T8338 = $signed(T8339) / $signed(22'h100000);
  assign T8339 = $signed(31'h3f174e6f) * $signed(16'h0);
  assign T8340 = {T8343, T8341};
  assign T8341 = $signed(T8342) / $signed(22'h100000);
  assign T8342 = $signed(29'h15407fbd) * $signed(16'h1);
  assign T8343 = T8344 ? 2'h3 : 2'h0;
  assign T8344 = T8341[6'h2c:6'h2c];
  assign T8345 = T2943[1'h0:1'h0];
  assign T8346 = T8361 ? twiddle4_3_191_real : twiddle4_3_190_real;
  assign twiddle4_3_190_real = T8349 + T8347;
  assign T8347 = $signed(T8348) / $signed(22'h100000);
  assign T8348 = $signed(31'h3efd4c53) * $signed(16'h0);
  assign T8349 = {T8352, T8350};
  assign T8350 = $signed(T8351) / $signed(22'h100000);
  assign T8351 = $signed(29'h14abf67e) * $signed(16'h1);
  assign T8352 = T8353 ? 2'h3 : 2'h0;
  assign T8353 = T8350[6'h2c:6'h2c];
  assign twiddle4_3_191_real = T8356 + T8354;
  assign T8354 = $signed(T8355) / $signed(22'h100000);
  assign T8355 = $signed(31'h3ee1ec86) * $signed(16'h0);
  assign T8356 = {T8359, T8357};
  assign T8357 = $signed(T8358) / $signed(22'h100000);
  assign T8358 = $signed(29'h1417ac23) * $signed(16'h1);
  assign T8359 = T8360 ? 2'h3 : 2'h0;
  assign T8360 = T8357[6'h2c:6'h2c];
  assign T8361 = T2943[1'h0:1'h0];
  assign T8362 = T2943[1'h1:1'h1];
  assign T8363 = T2943[2'h2:2'h2];
  assign T8364 = T2943[2'h3:2'h3];
  assign T8365 = T2943[3'h4:3'h4];
  assign T8366 = T2943[3'h5:3'h5];
  assign T8367 = T8827 ? T8629 : T8368;
  assign T8368 = T8628 ? T8502 : T8369;
  assign T8369 = T8501 ? T8439 : T8370;
  assign T8370 = T8438 ? T8405 : T8371;
  assign T8371 = T8404 ? T8388 : T8372;
  assign T8372 = T8387 ? twiddle4_3_193_real : twiddle4_3_192_real;
  assign twiddle4_3_192_real = T8375 + T8373;
  assign T8373 = $signed(T8374) / $signed(22'h100000);
  assign T8374 = $signed(31'h3ec52f9f) * $signed(16'h0);
  assign T8375 = {T8378, T8376};
  assign T8376 = $signed(T8377) / $signed(22'h100000);
  assign T8377 = $signed(29'h1383a3e2) * $signed(16'h1);
  assign T8378 = T8379 ? 2'h3 : 2'h0;
  assign T8379 = T8376[6'h2c:6'h2c];
  assign twiddle4_3_193_real = T8382 + T8380;
  assign T8380 = $signed(T8381) / $signed(22'h100000);
  assign T8381 = $signed(31'h3ea7163f) * $signed(16'h0);
  assign T8382 = {T8385, T8383};
  assign T8383 = $signed(T8384) / $signed(22'h100000);
  assign T8384 = $signed(29'h12efe0f3) * $signed(16'h1);
  assign T8385 = T8386 ? 2'h3 : 2'h0;
  assign T8386 = T8383[6'h2c:6'h2c];
  assign T8387 = T2943[1'h0:1'h0];
  assign T8388 = T8403 ? twiddle4_3_195_real : twiddle4_3_194_real;
  assign twiddle4_3_194_real = T8391 + T8389;
  assign T8389 = $signed(T8390) / $signed(22'h100000);
  assign T8390 = $signed(31'h3e87a10b) * $signed(16'h0);
  assign T8391 = {T8394, T8392};
  assign T8392 = $signed(T8393) / $signed(22'h100000);
  assign T8393 = $signed(29'h125c6689) * $signed(16'h1);
  assign T8394 = T8395 ? 2'h3 : 2'h0;
  assign T8395 = T8392[6'h2c:6'h2c];
  assign twiddle4_3_195_real = T8398 + T8396;
  assign T8396 = $signed(T8397) / $signed(22'h100000);
  assign T8397 = $signed(31'h3e66d0b4) * $signed(16'h0);
  assign T8398 = {T8401, T8399};
  assign T8399 = $signed(T8400) / $signed(22'h100000);
  assign T8400 = $signed(29'h11c937d7) * $signed(16'h1);
  assign T8401 = T8402 ? 2'h3 : 2'h0;
  assign T8402 = T8399[6'h2c:6'h2c];
  assign T8403 = T2943[1'h0:1'h0];
  assign T8404 = T2943[1'h1:1'h1];
  assign T8405 = T8437 ? T8422 : T8406;
  assign T8406 = T8421 ? twiddle4_3_197_real : twiddle4_3_196_real;
  assign twiddle4_3_196_real = T8409 + T8407;
  assign T8407 = $signed(T8408) / $signed(22'h100000);
  assign T8408 = $signed(31'h3e44a5ee) * $signed(16'h0);
  assign T8409 = {T8412, T8410};
  assign T8410 = $signed(T8411) / $signed(22'h100000);
  assign T8411 = $signed(29'h1136580e) * $signed(16'h1);
  assign T8412 = T8413 ? 2'h3 : 2'h0;
  assign T8413 = T8410[6'h2c:6'h2c];
  assign twiddle4_3_197_real = T8416 + T8414;
  assign T8414 = $signed(T8415) / $signed(22'h100000);
  assign T8415 = $signed(31'h3e212179) * $signed(16'h0);
  assign T8416 = {T8419, T8417};
  assign T8417 = $signed(T8418) / $signed(22'h100000);
  assign T8418 = $signed(29'h10a3ca5d) * $signed(16'h1);
  assign T8419 = T8420 ? 2'h3 : 2'h0;
  assign T8420 = T8417[6'h2c:6'h2c];
  assign T8421 = T2943[1'h0:1'h0];
  assign T8422 = T8436 ? twiddle4_3_199_real : twiddle4_3_198_real;
  assign twiddle4_3_198_real = T8425 + T8423;
  assign T8423 = $signed(T8424) / $signed(22'h100000);
  assign T8424 = $signed(31'h3dfc4418) * $signed(16'h0);
  assign T8425 = {T8428, T8426};
  assign T8426 = $signed(T8427) / $signed(22'h100000);
  assign T8427 = $signed(29'h101191f3) * $signed(16'h1);
  assign T8428 = T8429 ? 2'h3 : 2'h0;
  assign T8429 = T8426[6'h2c:6'h2c];
  assign twiddle4_3_199_real = T8432 + T8430;
  assign T8430 = $signed(T8431) / $signed(22'h100000);
  assign T8431 = $signed(31'h3dd60e98) * $signed(16'h0);
  assign T8432 = {T8435, T8433};
  assign T8433 = $signed(T8434) / $signed(22'h100000);
  assign T8434 = $signed(30'h2f7fb1fb) * $signed(16'h1);
  assign T8435 = T8433[6'h2d:6'h2d];
  assign T8436 = T2943[1'h0:1'h0];
  assign T8437 = T2943[1'h1:1'h1];
  assign T8438 = T2943[2'h2:2'h2];
  assign T8439 = T8500 ? T8470 : T8440;
  assign T8440 = T8469 ? T8455 : T8441;
  assign T8441 = T8454 ? twiddle4_3_201_real : twiddle4_3_200_real;
  assign twiddle4_3_200_real = T8444 + T8442;
  assign T8442 = $signed(T8443) / $signed(22'h100000);
  assign T8443 = $signed(31'h3dae81ce) * $signed(16'h0);
  assign T8444 = {T8447, T8445};
  assign T8445 = $signed(T8446) / $signed(22'h100000);
  assign T8446 = $signed(30'h2eee2d9e) * $signed(16'h1);
  assign T8447 = T8445[6'h2d:6'h2d];
  assign twiddle4_3_201_real = T8450 + T8448;
  assign T8448 = $signed(T8449) / $signed(22'h100000);
  assign T8449 = $signed(31'h3d859e96) * $signed(16'h0);
  assign T8450 = {T8453, T8451};
  assign T8451 = $signed(T8452) / $signed(22'h100000);
  assign T8452 = $signed(30'h2e5d0805) * $signed(16'h1);
  assign T8453 = T8451[6'h2d:6'h2d];
  assign T8454 = T2943[1'h0:1'h0];
  assign T8455 = T8468 ? twiddle4_3_203_real : twiddle4_3_202_real;
  assign twiddle4_3_202_real = T8458 + T8456;
  assign T8456 = $signed(T8457) / $signed(22'h100000);
  assign T8457 = $signed(31'h3d5b65d1) * $signed(16'h0);
  assign T8458 = {T8461, T8459};
  assign T8459 = $signed(T8460) / $signed(22'h100000);
  assign T8460 = $signed(30'h2dcc4455) * $signed(16'h1);
  assign T8461 = T8459[6'h2d:6'h2d];
  assign twiddle4_3_203_real = T8464 + T8462;
  assign T8462 = $signed(T8463) / $signed(22'h100000);
  assign T8463 = $signed(31'h3d2fd86c) * $signed(16'h0);
  assign T8464 = {T8467, T8465};
  assign T8465 = $signed(T8466) / $signed(22'h100000);
  assign T8466 = $signed(30'h2d3be5b2) * $signed(16'h1);
  assign T8467 = T8465[6'h2d:6'h2d];
  assign T8468 = T2943[1'h0:1'h0];
  assign T8469 = T2943[1'h1:1'h1];
  assign T8470 = T8499 ? T8485 : T8471;
  assign T8471 = T8484 ? twiddle4_3_205_real : twiddle4_3_204_real;
  assign twiddle4_3_204_real = T8474 + T8472;
  assign T8472 = $signed(T8473) / $signed(22'h100000);
  assign T8473 = $signed(31'h3d02f756) * $signed(16'h0);
  assign T8474 = {T8477, T8475};
  assign T8475 = $signed(T8476) / $signed(22'h100000);
  assign T8476 = $signed(30'h2cabef3e) * $signed(16'h1);
  assign T8477 = T8475[6'h2d:6'h2d];
  assign twiddle4_3_205_real = T8480 + T8478;
  assign T8478 = $signed(T8479) / $signed(22'h100000);
  assign T8479 = $signed(31'h3cd4c38a) * $signed(16'h0);
  assign T8480 = {T8483, T8481};
  assign T8481 = $signed(T8482) / $signed(22'h100000);
  assign T8482 = $signed(30'h2c1c6417) * $signed(16'h1);
  assign T8483 = T8481[6'h2d:6'h2d];
  assign T8484 = T2943[1'h0:1'h0];
  assign T8485 = T8498 ? twiddle4_3_207_real : twiddle4_3_206_real;
  assign twiddle4_3_206_real = T8488 + T8486;
  assign T8486 = $signed(T8487) / $signed(22'h100000);
  assign T8487 = $signed(31'h3ca53e08) * $signed(16'h0);
  assign T8488 = {T8491, T8489};
  assign T8489 = $signed(T8490) / $signed(22'h100000);
  assign T8490 = $signed(30'h2b8d475b) * $signed(16'h1);
  assign T8491 = T8489[6'h2d:6'h2d];
  assign twiddle4_3_207_real = T8494 + T8492;
  assign T8492 = $signed(T8493) / $signed(22'h100000);
  assign T8493 = $signed(31'h3c7467d8) * $signed(16'h0);
  assign T8494 = {T8497, T8495};
  assign T8495 = $signed(T8496) / $signed(22'h100000);
  assign T8496 = $signed(30'h2afe9c24) * $signed(16'h1);
  assign T8497 = T8495[6'h2d:6'h2d];
  assign T8498 = T2943[1'h0:1'h0];
  assign T8499 = T2943[1'h1:1'h1];
  assign T8500 = T2943[2'h2:2'h2];
  assign T8501 = T2943[2'h3:2'h3];
  assign T8502 = T8627 ? T8565 : T8503;
  assign T8503 = T8564 ? T8534 : T8504;
  assign T8504 = T8533 ? T8519 : T8505;
  assign T8505 = T8518 ? twiddle4_3_209_real : twiddle4_3_208_real;
  assign twiddle4_3_208_real = T8508 + T8506;
  assign T8506 = $signed(T8507) / $signed(22'h100000);
  assign T8507 = $signed(31'h3c424209) * $signed(16'h0);
  assign T8508 = {T8511, T8509};
  assign T8509 = $signed(T8510) / $signed(22'h100000);
  assign T8510 = $signed(30'h2a70658b) * $signed(16'h1);
  assign T8511 = T8509[6'h2d:6'h2d];
  assign twiddle4_3_209_real = T8514 + T8512;
  assign T8512 = $signed(T8513) / $signed(22'h100000);
  assign T8513 = $signed(31'h3c0ecdb2) * $signed(16'h0);
  assign T8514 = {T8517, T8515};
  assign T8515 = $signed(T8516) / $signed(22'h100000);
  assign T8516 = $signed(30'h29e2a6a4) * $signed(16'h1);
  assign T8517 = T8515[6'h2d:6'h2d];
  assign T8518 = T2943[1'h0:1'h0];
  assign T8519 = T8532 ? twiddle4_3_211_real : twiddle4_3_210_real;
  assign twiddle4_3_210_real = T8522 + T8520;
  assign T8520 = $signed(T8521) / $signed(22'h100000);
  assign T8521 = $signed(31'h3bda0bef) * $signed(16'h0);
  assign T8522 = {T8525, T8523};
  assign T8523 = $signed(T8524) / $signed(22'h100000);
  assign T8524 = $signed(30'h29556283) * $signed(16'h1);
  assign T8525 = T8523[6'h2d:6'h2d];
  assign twiddle4_3_211_real = T8528 + T8526;
  assign T8526 = $signed(T8527) / $signed(22'h100000);
  assign T8527 = $signed(31'h3ba3fde7) * $signed(16'h0);
  assign T8528 = {T8531, T8529};
  assign T8529 = $signed(T8530) / $signed(22'h100000);
  assign T8530 = $signed(30'h28c89c37) * $signed(16'h1);
  assign T8531 = T8529[6'h2d:6'h2d];
  assign T8532 = T2943[1'h0:1'h0];
  assign T8533 = T2943[1'h1:1'h1];
  assign T8534 = T8563 ? T8549 : T8535;
  assign T8535 = T8548 ? twiddle4_3_213_real : twiddle4_3_212_real;
  assign twiddle4_3_212_real = T8538 + T8536;
  assign T8536 = $signed(T8537) / $signed(22'h100000);
  assign T8537 = $signed(31'h3b6ca4c4) * $signed(16'h0);
  assign T8538 = {T8541, T8539};
  assign T8539 = $signed(T8540) / $signed(22'h100000);
  assign T8540 = $signed(30'h283c56cf) * $signed(16'h1);
  assign T8541 = T8539[6'h2d:6'h2d];
  assign twiddle4_3_213_real = T8544 + T8542;
  assign T8542 = $signed(T8543) / $signed(22'h100000);
  assign T8543 = $signed(31'h3b3401bb) * $signed(16'h0);
  assign T8544 = {T8547, T8545};
  assign T8545 = $signed(T8546) / $signed(22'h100000);
  assign T8546 = $signed(30'h27b09556) * $signed(16'h1);
  assign T8547 = T8545[6'h2d:6'h2d];
  assign T8548 = T2943[1'h0:1'h0];
  assign T8549 = T8562 ? twiddle4_3_215_real : twiddle4_3_214_real;
  assign twiddle4_3_214_real = T8552 + T8550;
  assign T8550 = $signed(T8551) / $signed(22'h100000);
  assign T8551 = $signed(31'h3afa1605) * $signed(16'h0);
  assign T8552 = {T8555, T8553};
  assign T8553 = $signed(T8554) / $signed(22'h100000);
  assign T8554 = $signed(30'h27255ad2) * $signed(16'h1);
  assign T8555 = T8553[6'h2d:6'h2d];
  assign twiddle4_3_215_real = T8558 + T8556;
  assign T8556 = $signed(T8557) / $signed(22'h100000);
  assign T8557 = $signed(31'h3abee2e5) * $signed(16'h0);
  assign T8558 = {T8561, T8559};
  assign T8559 = $signed(T8560) / $signed(22'h100000);
  assign T8560 = $signed(30'h269aaa49) * $signed(16'h1);
  assign T8561 = T8559[6'h2d:6'h2d];
  assign T8562 = T2943[1'h0:1'h0];
  assign T8563 = T2943[1'h1:1'h1];
  assign T8564 = T2943[2'h2:2'h2];
  assign T8565 = T8626 ? T8596 : T8566;
  assign T8566 = T8595 ? T8581 : T8567;
  assign T8567 = T8580 ? twiddle4_3_217_real : twiddle4_3_216_real;
  assign twiddle4_3_216_real = T8570 + T8568;
  assign T8568 = $signed(T8569) / $signed(22'h100000);
  assign T8569 = $signed(31'h3a8269a2) * $signed(16'h0);
  assign T8570 = {T8573, T8571};
  assign T8571 = $signed(T8572) / $signed(22'h100000);
  assign T8572 = $signed(30'h261086bd) * $signed(16'h1);
  assign T8573 = T8571[6'h2d:6'h2d];
  assign twiddle4_3_217_real = T8576 + T8574;
  assign T8574 = $signed(T8575) / $signed(22'h100000);
  assign T8575 = $signed(31'h3a44ab8d) * $signed(16'h0);
  assign T8576 = {T8579, T8577};
  assign T8577 = $signed(T8578) / $signed(22'h100000);
  assign T8578 = $signed(30'h2586f32d) * $signed(16'h1);
  assign T8579 = T8577[6'h2d:6'h2d];
  assign T8580 = T2943[1'h0:1'h0];
  assign T8581 = T8594 ? twiddle4_3_219_real : twiddle4_3_218_real;
  assign twiddle4_3_218_real = T8584 + T8582;
  assign T8582 = $signed(T8583) / $signed(22'h100000);
  assign T8583 = $signed(31'h3a05a9fd) * $signed(16'h0);
  assign T8584 = {T8587, T8585};
  assign T8585 = $signed(T8586) / $signed(22'h100000);
  assign T8586 = $signed(30'h24fdf294) * $signed(16'h1);
  assign T8587 = T8585[6'h2d:6'h2d];
  assign twiddle4_3_219_real = T8590 + T8588;
  assign T8588 = $signed(T8589) / $signed(22'h100000);
  assign T8589 = $signed(31'h39c5664f) * $signed(16'h0);
  assign T8590 = {T8593, T8591};
  assign T8591 = $signed(T8592) / $signed(22'h100000);
  assign T8592 = $signed(30'h247587ec) * $signed(16'h1);
  assign T8593 = T8591[6'h2d:6'h2d];
  assign T8594 = T2943[1'h0:1'h0];
  assign T8595 = T2943[1'h1:1'h1];
  assign T8596 = T8625 ? T8611 : T8597;
  assign T8597 = T8610 ? twiddle4_3_221_real : twiddle4_3_220_real;
  assign twiddle4_3_220_real = T8600 + T8598;
  assign T8598 = $signed(T8599) / $signed(22'h100000);
  assign T8599 = $signed(31'h3983e1e7) * $signed(16'h0);
  assign T8600 = {T8603, T8601};
  assign T8601 = $signed(T8602) / $signed(22'h100000);
  assign T8602 = $signed(30'h23edb628) * $signed(16'h1);
  assign T8603 = T8601[6'h2d:6'h2d];
  assign twiddle4_3_221_real = T8606 + T8604;
  assign T8604 = $signed(T8605) / $signed(22'h100000);
  assign T8605 = $signed(31'h39411e33) * $signed(16'h0);
  assign T8606 = {T8609, T8607};
  assign T8607 = $signed(T8608) / $signed(22'h100000);
  assign T8608 = $signed(30'h2366803d) * $signed(16'h1);
  assign T8609 = T8607[6'h2d:6'h2d];
  assign T8610 = T2943[1'h0:1'h0];
  assign T8611 = T8624 ? twiddle4_3_223_real : twiddle4_3_222_real;
  assign twiddle4_3_222_real = T8614 + T8612;
  assign T8612 = $signed(T8613) / $signed(22'h100000);
  assign T8613 = $signed(31'h38fd1ca4) * $signed(16'h0);
  assign T8614 = {T8617, T8615};
  assign T8615 = $signed(T8616) / $signed(22'h100000);
  assign T8616 = $signed(30'h22dfe918) * $signed(16'h1);
  assign T8617 = T8615[6'h2d:6'h2d];
  assign twiddle4_3_223_real = T8620 + T8618;
  assign T8618 = $signed(T8619) / $signed(22'h100000);
  assign T8619 = $signed(31'h38b7deb3) * $signed(16'h0);
  assign T8620 = {T8623, T8621};
  assign T8621 = $signed(T8622) / $signed(22'h100000);
  assign T8622 = $signed(30'h2259f3a4) * $signed(16'h1);
  assign T8623 = T8621[6'h2d:6'h2d];
  assign T8624 = T2943[1'h0:1'h0];
  assign T8625 = T2943[1'h1:1'h1];
  assign T8626 = T2943[2'h2:2'h2];
  assign T8627 = T2943[2'h3:2'h3];
  assign T8628 = T2943[3'h4:3'h4];
  assign T8629 = T8826 ? T8732 : T8630;
  assign T8630 = T8731 ? T8685 : T8631;
  assign T8631 = T8684 ? T8662 : T8632;
  assign T8632 = T8661 ? T8647 : T8633;
  assign T8633 = T8646 ? twiddle4_3_225_real : twiddle4_3_224_real;
  assign twiddle4_3_224_real = T8636 + T8634;
  assign T8634 = $signed(T8635) / $signed(22'h100000);
  assign T8635 = $signed(31'h387165e3) * $signed(16'h0);
  assign T8636 = {T8639, T8637};
  assign T8637 = $signed(T8638) / $signed(22'h100000);
  assign T8638 = $signed(30'h21d4a2c8) * $signed(16'h1);
  assign T8639 = T8637[6'h2d:6'h2d];
  assign twiddle4_3_225_real = T8642 + T8640;
  assign T8640 = $signed(T8641) / $signed(22'h100000);
  assign T8641 = $signed(31'h3829b3b8) * $signed(16'h0);
  assign T8642 = {T8645, T8643};
  assign T8643 = $signed(T8644) / $signed(22'h100000);
  assign T8644 = $signed(30'h214ff96b) * $signed(16'h1);
  assign T8645 = T8643[6'h2d:6'h2d];
  assign T8646 = T2943[1'h0:1'h0];
  assign T8647 = T8660 ? twiddle4_3_227_real : twiddle4_3_226_real;
  assign twiddle4_3_226_real = T8650 + T8648;
  assign T8648 = $signed(T8649) / $signed(22'h100000);
  assign T8649 = $signed(31'h37e0c9c2) * $signed(16'h0);
  assign T8650 = {T8653, T8651};
  assign T8651 = $signed(T8652) / $signed(22'h100000);
  assign T8652 = $signed(30'h20cbfa6a) * $signed(16'h1);
  assign T8653 = T8651[6'h2d:6'h2d];
  assign twiddle4_3_227_real = T8656 + T8654;
  assign T8654 = $signed(T8655) / $signed(22'h100000);
  assign T8655 = $signed(31'h3796a996) * $signed(16'h0);
  assign T8656 = {T8659, T8657};
  assign T8657 = $signed(T8658) / $signed(22'h100000);
  assign T8658 = $signed(30'h2048a8a4) * $signed(16'h1);
  assign T8659 = T8657[6'h2d:6'h2d];
  assign T8660 = T2943[1'h0:1'h0];
  assign T8661 = T2943[1'h1:1'h1];
  assign T8662 = T8683 ? T8673 : T8663;
  assign T8663 = T8672 ? twiddle4_3_229_real : twiddle4_3_228_real;
  assign twiddle4_3_228_real = T8666 + T8664;
  assign T8664 = $signed(T8665) / $signed(22'h100000);
  assign T8665 = $signed(31'h374b54ce) * $signed(16'h0);
  assign T8666 = $signed(T8667) / $signed(22'h100000);
  assign T8667 = $signed(31'h5fc606f2) * $signed(16'h1);
  assign twiddle4_3_229_real = T8670 + T8668;
  assign T8668 = $signed(T8669) / $signed(22'h100000);
  assign T8669 = $signed(31'h36fecd0d) * $signed(16'h0);
  assign T8670 = $signed(T8671) / $signed(22'h100000);
  assign T8671 = $signed(31'h5f441828) * $signed(16'h1);
  assign T8672 = T2943[1'h0:1'h0];
  assign T8673 = T8682 ? twiddle4_3_231_real : twiddle4_3_230_real;
  assign twiddle4_3_230_real = T8676 + T8674;
  assign T8674 = $signed(T8675) / $signed(22'h100000);
  assign T8675 = $signed(31'h36b113fd) * $signed(16'h0);
  assign T8676 = $signed(T8677) / $signed(22'h100000);
  assign T8677 = $signed(31'h5ec2df18) * $signed(16'h1);
  assign twiddle4_3_231_real = T8680 + T8678;
  assign T8678 = $signed(T8679) / $signed(22'h100000);
  assign T8679 = $signed(31'h36622b4b) * $signed(16'h0);
  assign T8680 = $signed(T8681) / $signed(22'h100000);
  assign T8681 = $signed(31'h5e425e90) * $signed(16'h1);
  assign T8682 = T2943[1'h0:1'h0];
  assign T8683 = T2943[1'h1:1'h1];
  assign T8684 = T2943[2'h2:2'h2];
  assign T8685 = T8730 ? T8708 : T8686;
  assign T8686 = T8707 ? T8697 : T8687;
  assign T8687 = T8696 ? twiddle4_3_233_real : twiddle4_3_232_real;
  assign twiddle4_3_232_real = T8690 + T8688;
  assign T8688 = $signed(T8689) / $signed(22'h100000);
  assign T8689 = $signed(31'h361214b0) * $signed(16'h0);
  assign T8690 = $signed(T8691) / $signed(22'h100000);
  assign T8691 = $signed(31'h5dc29958) * $signed(16'h1);
  assign twiddle4_3_233_real = T8694 + T8692;
  assign T8692 = $signed(T8693) / $signed(22'h100000);
  assign T8693 = $signed(31'h35c0d1e6) * $signed(16'h0);
  assign T8694 = $signed(T8695) / $signed(22'h100000);
  assign T8695 = $signed(31'h5d439237) * $signed(16'h1);
  assign T8696 = T2943[1'h0:1'h0];
  assign T8697 = T8706 ? twiddle4_3_235_real : twiddle4_3_234_real;
  assign twiddle4_3_234_real = T8700 + T8698;
  assign T8698 = $signed(T8699) / $signed(22'h100000);
  assign T8699 = $signed(31'h356e64b2) * $signed(16'h0);
  assign T8700 = $signed(T8701) / $signed(22'h100000);
  assign T8701 = $signed(31'h5cc54bed) * $signed(16'h1);
  assign twiddle4_3_235_real = T8704 + T8702;
  assign T8702 = $signed(T8703) / $signed(22'h100000);
  assign T8703 = $signed(31'h351acedc) * $signed(16'h0);
  assign T8704 = $signed(T8705) / $signed(22'h100000);
  assign T8705 = $signed(31'h5c47c937) * $signed(16'h1);
  assign T8706 = T2943[1'h0:1'h0];
  assign T8707 = T2943[1'h1:1'h1];
  assign T8708 = T8729 ? T8719 : T8709;
  assign T8709 = T8718 ? twiddle4_3_237_real : twiddle4_3_236_real;
  assign twiddle4_3_236_real = T8712 + T8710;
  assign T8710 = $signed(T8711) / $signed(22'h100000);
  assign T8711 = $signed(31'h34c61236) * $signed(16'h0);
  assign T8712 = $signed(T8713) / $signed(22'h100000);
  assign T8713 = $signed(31'h5bcb0cce) * $signed(16'h1);
  assign twiddle4_3_237_real = T8716 + T8714;
  assign T8714 = $signed(T8715) / $signed(22'h100000);
  assign T8715 = $signed(31'h34703094) * $signed(16'h0);
  assign T8716 = $signed(T8717) / $signed(22'h100000);
  assign T8717 = $signed(31'h5b4f1967) * $signed(16'h1);
  assign T8718 = T2943[1'h0:1'h0];
  assign T8719 = T8728 ? twiddle4_3_239_real : twiddle4_3_238_real;
  assign twiddle4_3_238_real = T8722 + T8720;
  assign T8720 = $signed(T8721) / $signed(22'h100000);
  assign T8721 = $signed(31'h34192bd5) * $signed(16'h0);
  assign T8722 = $signed(T8723) / $signed(22'h100000);
  assign T8723 = $signed(31'h5ad3f1b2) * $signed(16'h1);
  assign twiddle4_3_239_real = T8726 + T8724;
  assign T8724 = $signed(T8725) / $signed(22'h100000);
  assign T8725 = $signed(31'h33c105db) * $signed(16'h0);
  assign T8726 = $signed(T8727) / $signed(22'h100000);
  assign T8727 = $signed(31'h5a59985a) * $signed(16'h1);
  assign T8728 = T2943[1'h0:1'h0];
  assign T8729 = T2943[1'h1:1'h1];
  assign T8730 = T2943[2'h2:2'h2];
  assign T8731 = T2943[2'h3:2'h3];
  assign T8732 = T8825 ? T8779 : T8733;
  assign T8733 = T8778 ? T8756 : T8734;
  assign T8734 = T8755 ? T8745 : T8735;
  assign T8735 = T8744 ? twiddle4_3_241_real : twiddle4_3_240_real;
  assign twiddle4_3_240_real = T8738 + T8736;
  assign T8736 = $signed(T8737) / $signed(22'h100000);
  assign T8737 = $signed(31'h3367c08f) * $signed(16'h0);
  assign T8738 = $signed(T8739) / $signed(22'h100000);
  assign T8739 = $signed(31'h59e01007) * $signed(16'h1);
  assign twiddle4_3_241_real = T8742 + T8740;
  assign T8740 = $signed(T8741) / $signed(22'h100000);
  assign T8741 = $signed(31'h330d5de2) * $signed(16'h0);
  assign T8742 = $signed(T8743) / $signed(22'h100000);
  assign T8743 = $signed(31'h59675b5b) * $signed(16'h1);
  assign T8744 = T2943[1'h0:1'h0];
  assign T8745 = T8754 ? twiddle4_3_243_real : twiddle4_3_242_real;
  assign twiddle4_3_242_real = T8748 + T8746;
  assign T8746 = $signed(T8747) / $signed(22'h100000);
  assign T8747 = $signed(31'h32b1dfc9) * $signed(16'h0);
  assign T8748 = $signed(T8749) / $signed(22'h100000);
  assign T8749 = $signed(31'h58ef7cf5) * $signed(16'h1);
  assign twiddle4_3_243_real = T8752 + T8750;
  assign T8750 = $signed(T8751) / $signed(22'h100000);
  assign T8751 = $signed(31'h3255483f) * $signed(16'h0);
  assign T8752 = $signed(T8753) / $signed(22'h100000);
  assign T8753 = $signed(31'h5878776d) * $signed(16'h1);
  assign T8754 = T2943[1'h0:1'h0];
  assign T8755 = T2943[1'h1:1'h1];
  assign T8756 = T8777 ? T8767 : T8757;
  assign T8757 = T8766 ? twiddle4_3_245_real : twiddle4_3_244_real;
  assign twiddle4_3_244_real = T8760 + T8758;
  assign T8758 = $signed(T8759) / $signed(22'h100000);
  assign T8759 = $signed(31'h31f79947) * $signed(16'h0);
  assign T8760 = $signed(T8761) / $signed(22'h100000);
  assign T8761 = $signed(31'h58024d5a) * $signed(16'h1);
  assign twiddle4_3_245_real = T8764 + T8762;
  assign T8762 = $signed(T8763) / $signed(22'h100000);
  assign T8763 = $signed(31'h3198d4ea) * $signed(16'h0);
  assign T8764 = $signed(T8765) / $signed(22'h100000);
  assign T8765 = $signed(31'h578d014a) * $signed(16'h1);
  assign T8766 = T2943[1'h0:1'h0];
  assign T8767 = T8776 ? twiddle4_3_247_real : twiddle4_3_246_real;
  assign twiddle4_3_246_real = T8770 + T8768;
  assign T8768 = $signed(T8769) / $signed(22'h100000);
  assign T8769 = $signed(31'h3138fd34) * $signed(16'h0);
  assign T8770 = $signed(T8771) / $signed(22'h100000);
  assign T8771 = $signed(31'h571895c9) * $signed(16'h1);
  assign twiddle4_3_247_real = T8774 + T8772;
  assign T8772 = $signed(T8773) / $signed(22'h100000);
  assign T8773 = $signed(31'h30d8143b) * $signed(16'h0);
  assign T8774 = $signed(T8775) / $signed(22'h100000);
  assign T8775 = $signed(31'h56a50d5e) * $signed(16'h1);
  assign T8776 = T2943[1'h0:1'h0];
  assign T8777 = T2943[1'h1:1'h1];
  assign T8778 = T2943[2'h2:2'h2];
  assign T8779 = T8824 ? T8802 : T8780;
  assign T8780 = T8801 ? T8791 : T8781;
  assign T8781 = T8790 ? twiddle4_3_249_real : twiddle4_3_248_real;
  assign twiddle4_3_248_real = T8784 + T8782;
  assign T8782 = $signed(T8783) / $signed(22'h100000);
  assign T8783 = $signed(31'h30761c17) * $signed(16'h0);
  assign T8784 = $signed(T8785) / $signed(22'h100000);
  assign T8785 = $signed(31'h56326a89) * $signed(16'h1);
  assign twiddle4_3_249_real = T8788 + T8786;
  assign T8786 = $signed(T8787) / $signed(22'h100000);
  assign T8787 = $signed(31'h301316ea) * $signed(16'h0);
  assign T8788 = $signed(T8789) / $signed(22'h100000);
  assign T8789 = $signed(31'h55c0afc7) * $signed(16'h1);
  assign T8790 = T2943[1'h0:1'h0];
  assign T8791 = T8800 ? twiddle4_3_251_real : twiddle4_3_250_real;
  assign twiddle4_3_250_real = T8794 + T8792;
  assign T8792 = $signed(T8793) / $signed(22'h100000);
  assign T8793 = $signed(31'h2faf06d9) * $signed(16'h0);
  assign T8794 = $signed(T8795) / $signed(22'h100000);
  assign T8795 = $signed(31'h554fdf8f) * $signed(16'h1);
  assign twiddle4_3_251_real = T8798 + T8796;
  assign T8796 = $signed(T8797) / $signed(22'h100000);
  assign T8797 = $signed(31'h2f49ee0f) * $signed(16'h0);
  assign T8798 = $signed(T8799) / $signed(22'h100000);
  assign T8799 = $signed(31'h54dffc55) * $signed(16'h1);
  assign T8800 = T2943[1'h0:1'h0];
  assign T8801 = T2943[1'h1:1'h1];
  assign T8802 = T8823 ? T8813 : T8803;
  assign T8803 = T8812 ? twiddle4_3_253_real : twiddle4_3_252_real;
  assign twiddle4_3_252_real = T8806 + T8804;
  assign T8804 = $signed(T8805) / $signed(22'h100000);
  assign T8805 = $signed(31'h2ee3cebe) * $signed(16'h0);
  assign T8806 = $signed(T8807) / $signed(22'h100000);
  assign T8807 = $signed(31'h54710884) * $signed(16'h1);
  assign twiddle4_3_253_real = T8810 + T8808;
  assign T8808 = $signed(T8809) / $signed(22'h100000);
  assign T8809 = $signed(31'h2e7cab1c) * $signed(16'h0);
  assign T8810 = $signed(T8811) / $signed(22'h100000);
  assign T8811 = $signed(31'h54030685) * $signed(16'h1);
  assign T8812 = T2943[1'h0:1'h0];
  assign T8813 = T8822 ? twiddle4_3_255_real : twiddle4_3_254_real;
  assign twiddle4_3_254_real = T8816 + T8814;
  assign T8814 = $signed(T8815) / $signed(22'h100000);
  assign T8815 = $signed(31'h2e148566) * $signed(16'h0);
  assign T8816 = $signed(T8817) / $signed(22'h100000);
  assign T8817 = $signed(31'h5395f8ba) * $signed(16'h1);
  assign twiddle4_3_255_real = T8820 + T8818;
  assign T8818 = $signed(T8819) / $signed(22'h100000);
  assign T8819 = $signed(31'h2dab5fde) * $signed(16'h0);
  assign T8820 = $signed(T8821) / $signed(22'h100000);
  assign T8821 = $signed(31'h5329e182) * $signed(16'h1);
  assign T8822 = T2943[1'h0:1'h0];
  assign T8823 = T2943[1'h1:1'h1];
  assign T8824 = T2943[2'h2:2'h2];
  assign T8825 = T2943[2'h3:2'h3];
  assign T8826 = T2943[3'h4:3'h4];
  assign T8827 = T2943[3'h5:3'h5];
  assign T8828 = T2943[3'h6:3'h6];
  assign T8829 = T7808[6'h2e:6'h2e];
  assign T8830 = T2943[3'h7:3'h7];
  assign T8831 = {T10788, T8832};
  assign T8832 = T10787 ? T9852 : T8833;
  assign T8833 = T9851 ? T9292 : T8834;
  assign T8834 = T9291 ? T9031 : T8835;
  assign T8835 = T9030 ? T8930 : T8836;
  assign T8836 = T8929 ? T8883 : T8837;
  assign T8837 = T8882 ? T8860 : T8838;
  assign T8838 = T8859 ? T8849 : T8839;
  assign T8839 = T8848 ? twiddle4_3_257_real : twiddle4_3_256_real;
  assign twiddle4_3_256_real = T8842 + T8840;
  assign T8840 = $signed(T8841) / $signed(22'h100000);
  assign T8841 = $signed(31'h2d413ccc) * $signed(16'h0);
  assign T8842 = $signed(T8843) / $signed(22'h100000);
  assign T8843 = $signed(31'h52bec334) * $signed(16'h1);
  assign twiddle4_3_257_real = T8846 + T8844;
  assign T8844 = $signed(T8845) / $signed(22'h100000);
  assign T8845 = $signed(31'h2cd61e7e) * $signed(16'h0);
  assign T8846 = $signed(T8847) / $signed(22'h100000);
  assign T8847 = $signed(31'h5254a022) * $signed(16'h1);
  assign T8848 = T2943[1'h0:1'h0];
  assign T8849 = T8858 ? twiddle4_3_259_real : twiddle4_3_258_real;
  assign twiddle4_3_258_real = T8852 + T8850;
  assign T8850 = $signed(T8851) / $signed(22'h100000);
  assign T8851 = $signed(31'h2c6a0746) * $signed(16'h0);
  assign T8852 = $signed(T8853) / $signed(22'h100000);
  assign T8853 = $signed(31'h51eb7a9a) * $signed(16'h1);
  assign twiddle4_3_259_real = T8856 + T8854;
  assign T8854 = $signed(T8855) / $signed(22'h100000);
  assign T8855 = $signed(31'h2bfcf97b) * $signed(16'h0);
  assign T8856 = $signed(T8857) / $signed(22'h100000);
  assign T8857 = $signed(31'h518354e4) * $signed(16'h1);
  assign T8858 = T2943[1'h0:1'h0];
  assign T8859 = T2943[1'h1:1'h1];
  assign T8860 = T8881 ? T8871 : T8861;
  assign T8861 = T8870 ? twiddle4_3_261_real : twiddle4_3_260_real;
  assign twiddle4_3_260_real = T8864 + T8862;
  assign T8862 = $signed(T8863) / $signed(22'h100000);
  assign T8863 = $signed(31'h2b8ef77c) * $signed(16'h0);
  assign T8864 = $signed(T8865) / $signed(22'h100000);
  assign T8865 = $signed(31'h511c3142) * $signed(16'h1);
  assign twiddle4_3_261_real = T8868 + T8866;
  assign T8866 = $signed(T8867) / $signed(22'h100000);
  assign T8867 = $signed(31'h2b2003ab) * $signed(16'h0);
  assign T8868 = $signed(T8869) / $signed(22'h100000);
  assign T8869 = $signed(31'h50b611f1) * $signed(16'h1);
  assign T8870 = T2943[1'h0:1'h0];
  assign T8871 = T8880 ? twiddle4_3_263_real : twiddle4_3_262_real;
  assign twiddle4_3_262_real = T8874 + T8872;
  assign T8872 = $signed(T8873) / $signed(22'h100000);
  assign T8873 = $signed(31'h2ab02071) * $signed(16'h0);
  assign T8874 = $signed(T8875) / $signed(22'h100000);
  assign T8875 = $signed(31'h5050f927) * $signed(16'h1);
  assign twiddle4_3_263_real = T8878 + T8876;
  assign T8876 = $signed(T8877) / $signed(22'h100000);
  assign T8877 = $signed(31'h2a3f5039) * $signed(16'h0);
  assign T8878 = $signed(T8879) / $signed(22'h100000);
  assign T8879 = $signed(31'h4fece916) * $signed(16'h1);
  assign T8880 = T2943[1'h0:1'h0];
  assign T8881 = T2943[1'h1:1'h1];
  assign T8882 = T2943[2'h2:2'h2];
  assign T8883 = T8928 ? T8906 : T8884;
  assign T8884 = T8905 ? T8895 : T8885;
  assign T8885 = T8894 ? twiddle4_3_265_real : twiddle4_3_264_real;
  assign twiddle4_3_264_real = T8888 + T8886;
  assign T8886 = $signed(T8887) / $signed(22'h100000);
  assign T8887 = $signed(31'h29cd9577) * $signed(16'h0);
  assign T8888 = $signed(T8889) / $signed(22'h100000);
  assign T8889 = $signed(31'h4f89e3e9) * $signed(16'h1);
  assign twiddle4_3_265_real = T8892 + T8890;
  assign T8890 = $signed(T8891) / $signed(22'h100000);
  assign T8891 = $signed(31'h295af2a2) * $signed(16'h0);
  assign T8892 = $signed(T8893) / $signed(22'h100000);
  assign T8893 = $signed(31'h4f27ebc5) * $signed(16'h1);
  assign T8894 = T2943[1'h0:1'h0];
  assign T8895 = T8904 ? twiddle4_3_267_real : twiddle4_3_266_real;
  assign twiddle4_3_266_real = T8898 + T8896;
  assign T8896 = $signed(T8897) / $signed(22'h100000);
  assign T8897 = $signed(31'h28e76a37) * $signed(16'h0);
  assign T8898 = $signed(T8899) / $signed(22'h100000);
  assign T8899 = $signed(31'h4ec702cc) * $signed(16'h1);
  assign twiddle4_3_267_real = T8902 + T8900;
  assign T8900 = $signed(T8901) / $signed(22'h100000);
  assign T8901 = $signed(31'h2872feb6) * $signed(16'h0);
  assign T8902 = $signed(T8903) / $signed(22'h100000);
  assign T8903 = $signed(31'h4e672b16) * $signed(16'h1);
  assign T8904 = T2943[1'h0:1'h0];
  assign T8905 = T2943[1'h1:1'h1];
  assign T8906 = T8927 ? T8917 : T8907;
  assign T8907 = T8916 ? twiddle4_3_269_real : twiddle4_3_268_real;
  assign twiddle4_3_268_real = T8910 + T8908;
  assign T8908 = $signed(T8909) / $signed(22'h100000);
  assign T8909 = $signed(31'h27fdb2a6) * $signed(16'h0);
  assign T8910 = $signed(T8911) / $signed(22'h100000);
  assign T8911 = $signed(31'h4e0866b9) * $signed(16'h1);
  assign twiddle4_3_269_real = T8914 + T8912;
  assign T8912 = $signed(T8913) / $signed(22'h100000);
  assign T8913 = $signed(31'h27878893) * $signed(16'h0);
  assign T8914 = $signed(T8915) / $signed(22'h100000);
  assign T8915 = $signed(31'h4daab7c1) * $signed(16'h1);
  assign T8916 = T2943[1'h0:1'h0];
  assign T8917 = T8926 ? twiddle4_3_271_real : twiddle4_3_270_real;
  assign twiddle4_3_270_real = T8920 + T8918;
  assign T8918 = $signed(T8919) / $signed(22'h100000);
  assign T8919 = $signed(31'h2710830b) * $signed(16'h0);
  assign T8920 = $signed(T8921) / $signed(22'h100000);
  assign T8921 = $signed(31'h4d4e2037) * $signed(16'h1);
  assign twiddle4_3_271_real = T8924 + T8922;
  assign T8922 = $signed(T8923) / $signed(22'h100000);
  assign T8923 = $signed(31'h2698a4a5) * $signed(16'h0);
  assign T8924 = $signed(T8925) / $signed(22'h100000);
  assign T8925 = $signed(31'h4cf2a21e) * $signed(16'h1);
  assign T8926 = T2943[1'h0:1'h0];
  assign T8927 = T2943[1'h1:1'h1];
  assign T8928 = T2943[2'h2:2'h2];
  assign T8929 = T2943[2'h3:2'h3];
  assign T8930 = T9029 ? T8977 : T8931;
  assign T8931 = T8976 ? T8954 : T8932;
  assign T8932 = T8953 ? T8943 : T8933;
  assign T8933 = T8942 ? twiddle4_3_273_real : twiddle4_3_272_real;
  assign twiddle4_3_272_real = T8936 + T8934;
  assign T8934 = $signed(T8935) / $signed(22'h100000);
  assign T8935 = $signed(31'h261feff9) * $signed(16'h0);
  assign T8936 = $signed(T8937) / $signed(22'h100000);
  assign T8937 = $signed(31'h4c983f71) * $signed(16'h1);
  assign twiddle4_3_273_real = T8940 + T8938;
  assign T8938 = $signed(T8939) / $signed(22'h100000);
  assign T8939 = $signed(31'h25a667a6) * $signed(16'h0);
  assign T8940 = $signed(T8941) / $signed(22'h100000);
  assign T8941 = $signed(31'h4c3efa25) * $signed(16'h1);
  assign T8942 = T2943[1'h0:1'h0];
  assign T8943 = T8952 ? twiddle4_3_275_real : twiddle4_3_274_real;
  assign twiddle4_3_274_real = T8946 + T8944;
  assign T8944 = $signed(T8945) / $signed(22'h100000);
  assign T8945 = $signed(31'h252c0e4e) * $signed(16'h0);
  assign T8946 = $signed(T8947) / $signed(22'h100000);
  assign T8947 = $signed(31'h4be6d42b) * $signed(16'h1);
  assign twiddle4_3_275_real = T8950 + T8948;
  assign T8948 = $signed(T8949) / $signed(22'h100000);
  assign T8949 = $signed(31'h24b0e699) * $signed(16'h0);
  assign T8950 = $signed(T8951) / $signed(22'h100000);
  assign T8951 = $signed(31'h4b8fcf6c) * $signed(16'h1);
  assign T8952 = T2943[1'h0:1'h0];
  assign T8953 = T2943[1'h1:1'h1];
  assign T8954 = T8975 ? T8965 : T8955;
  assign T8955 = T8964 ? twiddle4_3_277_real : twiddle4_3_276_real;
  assign twiddle4_3_276_real = T8958 + T8956;
  assign T8956 = $signed(T8957) / $signed(22'h100000);
  assign T8957 = $signed(31'h2434f332) * $signed(16'h0);
  assign T8958 = $signed(T8959) / $signed(22'h100000);
  assign T8959 = $signed(31'h4b39edca) * $signed(16'h1);
  assign twiddle4_3_277_real = T8962 + T8960;
  assign T8960 = $signed(T8961) / $signed(22'h100000);
  assign T8961 = $signed(31'h23b836c9) * $signed(16'h0);
  assign T8962 = $signed(T8963) / $signed(22'h100000);
  assign T8963 = $signed(31'h4ae53124) * $signed(16'h1);
  assign T8964 = T2943[1'h0:1'h0];
  assign T8965 = T8974 ? twiddle4_3_279_real : twiddle4_3_278_real;
  assign twiddle4_3_278_real = T8968 + T8966;
  assign T8966 = $signed(T8967) / $signed(22'h100000);
  assign T8967 = $signed(31'h233ab413) * $signed(16'h0);
  assign T8968 = $signed(T8969) / $signed(22'h100000);
  assign T8969 = $signed(31'h4a919b4e) * $signed(16'h1);
  assign twiddle4_3_279_real = T8972 + T8970;
  assign T8970 = $signed(T8971) / $signed(22'h100000);
  assign T8971 = $signed(31'h22bc6dc9) * $signed(16'h0);
  assign T8972 = $signed(T8973) / $signed(22'h100000);
  assign T8973 = $signed(31'h4a3f2e1a) * $signed(16'h1);
  assign T8974 = T2943[1'h0:1'h0];
  assign T8975 = T2943[1'h1:1'h1];
  assign T8976 = T2943[2'h2:2'h2];
  assign T8977 = T9028 ? T9000 : T8978;
  assign T8978 = T8999 ? T8989 : T8979;
  assign T8979 = T8988 ? twiddle4_3_281_real : twiddle4_3_280_real;
  assign twiddle4_3_280_real = T8982 + T8980;
  assign T8980 = $signed(T8981) / $signed(22'h100000);
  assign T8981 = $signed(31'h223d66a8) * $signed(16'h0);
  assign T8982 = $signed(T8983) / $signed(22'h100000);
  assign T8983 = $signed(31'h49edeb50) * $signed(16'h1);
  assign twiddle4_3_281_real = T8986 + T8984;
  assign T8984 = $signed(T8985) / $signed(22'h100000);
  assign T8985 = $signed(31'h21bda170) * $signed(16'h0);
  assign T8986 = $signed(T8987) / $signed(22'h100000);
  assign T8987 = $signed(31'h499dd4b5) * $signed(16'h1);
  assign T8988 = T2943[1'h0:1'h0];
  assign T8989 = T8998 ? twiddle4_3_283_real : twiddle4_3_282_real;
  assign twiddle4_3_282_real = T8992 + T8990;
  assign T8990 = $signed(T8991) / $signed(22'h100000);
  assign T8991 = $signed(31'h213d20e8) * $signed(16'h0);
  assign T8992 = $signed(T8993) / $signed(22'h100000);
  assign T8993 = $signed(31'h494eec03) * $signed(16'h1);
  assign twiddle4_3_283_real = T8996 + T8994;
  assign T8994 = $signed(T8995) / $signed(22'h100000);
  assign T8995 = $signed(31'h20bbe7d8) * $signed(16'h0);
  assign T8996 = $signed(T8997) / $signed(22'h100000);
  assign T8997 = $signed(31'h490132f3) * $signed(16'h1);
  assign T8998 = T2943[1'h0:1'h0];
  assign T8999 = T2943[1'h1:1'h1];
  assign T9000 = T9027 ? T9013 : T9001;
  assign T9001 = T9012 ? twiddle4_3_285_real : twiddle4_3_284_real;
  assign twiddle4_3_284_real = T9004 + T9002;
  assign T9002 = $signed(T9003) / $signed(22'h100000);
  assign T9003 = $signed(31'h2039f90e) * $signed(16'h0);
  assign T9004 = $signed(T9005) / $signed(22'h100000);
  assign T9005 = $signed(31'h48b4ab32) * $signed(16'h1);
  assign twiddle4_3_285_real = T9010 + T9006;
  assign T9006 = {T9009, T9007};
  assign T9007 = $signed(T9008) / $signed(22'h100000);
  assign T9008 = $signed(30'h1fb7575c) * $signed(16'h0);
  assign T9009 = T9007[6'h2d:6'h2d];
  assign T9010 = $signed(T9011) / $signed(22'h100000);
  assign T9011 = $signed(31'h4869566a) * $signed(16'h1);
  assign T9012 = T2943[1'h0:1'h0];
  assign T9013 = T9026 ? twiddle4_3_287_real : twiddle4_3_286_real;
  assign twiddle4_3_286_real = T9018 + T9014;
  assign T9014 = {T9017, T9015};
  assign T9015 = $signed(T9016) / $signed(22'h100000);
  assign T9016 = $signed(30'h1f340596) * $signed(16'h0);
  assign T9017 = T9015[6'h2d:6'h2d];
  assign T9018 = $signed(T9019) / $signed(22'h100000);
  assign T9019 = $signed(31'h481f363e) * $signed(16'h1);
  assign twiddle4_3_287_real = T9024 + T9020;
  assign T9020 = {T9023, T9021};
  assign T9021 = $signed(T9022) / $signed(22'h100000);
  assign T9022 = $signed(30'h1eb00695) * $signed(16'h0);
  assign T9023 = T9021[6'h2d:6'h2d];
  assign T9024 = $signed(T9025) / $signed(22'h100000);
  assign T9025 = $signed(31'h47d64c48) * $signed(16'h1);
  assign T9026 = T2943[1'h0:1'h0];
  assign T9027 = T2943[1'h1:1'h1];
  assign T9028 = T2943[2'h2:2'h2];
  assign T9029 = T2943[2'h3:2'h3];
  assign T9030 = T2943[3'h4:3'h4];
  assign T9031 = T9290 ? T9158 : T9032;
  assign T9032 = T9157 ? T9095 : T9033;
  assign T9033 = T9094 ? T9064 : T9034;
  assign T9034 = T9063 ? T9049 : T9035;
  assign T9035 = T9048 ? twiddle4_3_289_real : twiddle4_3_288_real;
  assign twiddle4_3_288_real = T9040 + T9036;
  assign T9036 = {T9039, T9037};
  assign T9037 = $signed(T9038) / $signed(22'h100000);
  assign T9038 = $signed(30'h1e2b5d38) * $signed(16'h0);
  assign T9039 = T9037[6'h2d:6'h2d];
  assign T9040 = $signed(T9041) / $signed(22'h100000);
  assign T9041 = $signed(31'h478e9a1d) * $signed(16'h1);
  assign twiddle4_3_289_real = T9046 + T9042;
  assign T9042 = {T9045, T9043};
  assign T9043 = $signed(T9044) / $signed(22'h100000);
  assign T9044 = $signed(30'h1da60c5c) * $signed(16'h0);
  assign T9045 = T9043[6'h2d:6'h2d];
  assign T9046 = $signed(T9047) / $signed(22'h100000);
  assign T9047 = $signed(31'h4748214d) * $signed(16'h1);
  assign T9048 = T2943[1'h0:1'h0];
  assign T9049 = T9062 ? twiddle4_3_291_real : twiddle4_3_290_real;
  assign twiddle4_3_290_real = T9054 + T9050;
  assign T9050 = {T9053, T9051};
  assign T9051 = $signed(T9052) / $signed(22'h100000);
  assign T9052 = $signed(30'h1d2016e8) * $signed(16'h0);
  assign T9053 = T9051[6'h2d:6'h2d];
  assign T9054 = $signed(T9055) / $signed(22'h100000);
  assign T9055 = $signed(31'h4702e35c) * $signed(16'h1);
  assign twiddle4_3_291_real = T9060 + T9056;
  assign T9056 = {T9059, T9057};
  assign T9057 = $signed(T9058) / $signed(22'h100000);
  assign T9058 = $signed(30'h1c997fc3) * $signed(16'h0);
  assign T9059 = T9057[6'h2d:6'h2d];
  assign T9060 = $signed(T9061) / $signed(22'h100000);
  assign T9061 = $signed(31'h46bee1cd) * $signed(16'h1);
  assign T9062 = T2943[1'h0:1'h0];
  assign T9063 = T2943[1'h1:1'h1];
  assign T9064 = T9093 ? T9079 : T9065;
  assign T9065 = T9078 ? twiddle4_3_293_real : twiddle4_3_292_real;
  assign twiddle4_3_292_real = T9070 + T9066;
  assign T9066 = {T9069, T9067};
  assign T9067 = $signed(T9068) / $signed(22'h100000);
  assign T9068 = $signed(30'h1c1249d8) * $signed(16'h0);
  assign T9069 = T9067[6'h2d:6'h2d];
  assign T9070 = $signed(T9071) / $signed(22'h100000);
  assign T9071 = $signed(31'h467c1e19) * $signed(16'h1);
  assign twiddle4_3_293_real = T9076 + T9072;
  assign T9072 = {T9075, T9073};
  assign T9073 = $signed(T9074) / $signed(22'h100000);
  assign T9074 = $signed(30'h1b8a7814) * $signed(16'h0);
  assign T9075 = T9073[6'h2d:6'h2d];
  assign T9076 = $signed(T9077) / $signed(22'h100000);
  assign T9077 = $signed(31'h463a99b1) * $signed(16'h1);
  assign T9078 = T2943[1'h0:1'h0];
  assign T9079 = T9092 ? twiddle4_3_295_real : twiddle4_3_294_real;
  assign twiddle4_3_294_real = T9084 + T9080;
  assign T9080 = {T9083, T9081};
  assign T9081 = $signed(T9082) / $signed(22'h100000);
  assign T9082 = $signed(30'h1b020d6c) * $signed(16'h0);
  assign T9083 = T9081[6'h2d:6'h2d];
  assign T9084 = $signed(T9085) / $signed(22'h100000);
  assign T9085 = $signed(31'h45fa5603) * $signed(16'h1);
  assign twiddle4_3_295_real = T9090 + T9086;
  assign T9086 = {T9089, T9087};
  assign T9087 = $signed(T9088) / $signed(22'h100000);
  assign T9088 = $signed(30'h1a790cd3) * $signed(16'h0);
  assign T9089 = T9087[6'h2d:6'h2d];
  assign T9090 = $signed(T9091) / $signed(22'h100000);
  assign T9091 = $signed(31'h45bb5473) * $signed(16'h1);
  assign T9092 = T2943[1'h0:1'h0];
  assign T9093 = T2943[1'h1:1'h1];
  assign T9094 = T2943[2'h2:2'h2];
  assign T9095 = T9156 ? T9126 : T9096;
  assign T9096 = T9125 ? T9111 : T9097;
  assign T9097 = T9110 ? twiddle4_3_297_real : twiddle4_3_296_real;
  assign twiddle4_3_296_real = T9102 + T9098;
  assign T9098 = {T9101, T9099};
  assign T9099 = $signed(T9100) / $signed(22'h100000);
  assign T9100 = $signed(30'h19ef7943) * $signed(16'h0);
  assign T9101 = T9099[6'h2d:6'h2d];
  assign T9102 = $signed(T9103) / $signed(22'h100000);
  assign T9103 = $signed(31'h457d965e) * $signed(16'h1);
  assign twiddle4_3_297_real = T9108 + T9104;
  assign T9104 = {T9107, T9105};
  assign T9105 = $signed(T9106) / $signed(22'h100000);
  assign T9106 = $signed(30'h196555b7) * $signed(16'h0);
  assign T9107 = T9105[6'h2d:6'h2d];
  assign T9108 = $signed(T9109) / $signed(22'h100000);
  assign T9109 = $signed(31'h45411d1b) * $signed(16'h1);
  assign T9110 = T2943[1'h0:1'h0];
  assign T9111 = T9124 ? twiddle4_3_299_real : twiddle4_3_298_real;
  assign twiddle4_3_298_real = T9116 + T9112;
  assign T9112 = {T9115, T9113};
  assign T9113 = $signed(T9114) / $signed(22'h100000);
  assign T9114 = $signed(30'h18daa52e) * $signed(16'h0);
  assign T9115 = T9113[6'h2d:6'h2d];
  assign T9116 = $signed(T9117) / $signed(22'h100000);
  assign T9117 = $signed(31'h4505e9fb) * $signed(16'h1);
  assign twiddle4_3_299_real = T9122 + T9118;
  assign T9118 = {T9121, T9119};
  assign T9119 = $signed(T9120) / $signed(22'h100000);
  assign T9120 = $signed(30'h184f6aaa) * $signed(16'h0);
  assign T9121 = T9119[6'h2d:6'h2d];
  assign T9122 = $signed(T9123) / $signed(22'h100000);
  assign T9123 = $signed(31'h44cbfe45) * $signed(16'h1);
  assign T9124 = T2943[1'h0:1'h0];
  assign T9125 = T2943[1'h1:1'h1];
  assign T9126 = T9155 ? T9141 : T9127;
  assign T9127 = T9140 ? twiddle4_3_301_real : twiddle4_3_300_real;
  assign twiddle4_3_300_real = T9132 + T9128;
  assign T9128 = {T9131, T9129};
  assign T9129 = $signed(T9130) / $signed(22'h100000);
  assign T9130 = $signed(30'h17c3a931) * $signed(16'h0);
  assign T9131 = T9129[6'h2d:6'h2d];
  assign T9132 = $signed(T9133) / $signed(22'h100000);
  assign T9133 = $signed(31'h44935b3c) * $signed(16'h1);
  assign twiddle4_3_301_real = T9138 + T9134;
  assign T9134 = {T9137, T9135};
  assign T9135 = $signed(T9136) / $signed(22'h100000);
  assign T9136 = $signed(30'h173763c9) * $signed(16'h0);
  assign T9137 = T9135[6'h2d:6'h2d];
  assign T9138 = $signed(T9139) / $signed(22'h100000);
  assign T9139 = $signed(31'h445c0219) * $signed(16'h1);
  assign T9140 = T2943[1'h0:1'h0];
  assign T9141 = T9154 ? twiddle4_3_303_real : twiddle4_3_302_real;
  assign twiddle4_3_302_real = T9146 + T9142;
  assign T9142 = {T9145, T9143};
  assign T9143 = $signed(T9144) / $signed(22'h100000);
  assign T9144 = $signed(30'h16aa9d7d) * $signed(16'h0);
  assign T9145 = T9143[6'h2d:6'h2d];
  assign T9146 = $signed(T9147) / $signed(22'h100000);
  assign T9147 = $signed(31'h4425f411) * $signed(16'h1);
  assign twiddle4_3_303_real = T9152 + T9148;
  assign T9148 = {T9151, T9149};
  assign T9149 = $signed(T9150) / $signed(22'h100000);
  assign T9150 = $signed(30'h161d595c) * $signed(16'h0);
  assign T9151 = T9149[6'h2d:6'h2d];
  assign T9152 = $signed(T9153) / $signed(22'h100000);
  assign T9153 = $signed(31'h43f1324e) * $signed(16'h1);
  assign T9154 = T2943[1'h0:1'h0];
  assign T9155 = T2943[1'h1:1'h1];
  assign T9156 = T2943[2'h2:2'h2];
  assign T9157 = T2943[2'h3:2'h3];
  assign T9158 = T9289 ? T9221 : T9159;
  assign T9159 = T9220 ? T9190 : T9160;
  assign T9160 = T9189 ? T9175 : T9161;
  assign T9161 = T9174 ? twiddle4_3_305_real : twiddle4_3_304_real;
  assign twiddle4_3_304_real = T9166 + T9162;
  assign T9162 = {T9165, T9163};
  assign T9163 = $signed(T9164) / $signed(22'h100000);
  assign T9164 = $signed(30'h158f9a75) * $signed(16'h0);
  assign T9165 = T9163[6'h2d:6'h2d];
  assign T9166 = $signed(T9167) / $signed(22'h100000);
  assign T9167 = $signed(31'h43bdbdf7) * $signed(16'h1);
  assign twiddle4_3_305_real = T9172 + T9168;
  assign T9168 = {T9171, T9169};
  assign T9169 = $signed(T9170) / $signed(22'h100000);
  assign T9170 = $signed(30'h150163dc) * $signed(16'h0);
  assign T9171 = T9169[6'h2d:6'h2d];
  assign T9172 = $signed(T9173) / $signed(22'h100000);
  assign T9173 = $signed(31'h438b9828) * $signed(16'h1);
  assign T9174 = T2943[1'h0:1'h0];
  assign T9175 = T9188 ? twiddle4_3_307_real : twiddle4_3_306_real;
  assign twiddle4_3_306_real = T9180 + T9176;
  assign T9176 = {T9179, T9177};
  assign T9177 = $signed(T9178) / $signed(22'h100000);
  assign T9178 = $signed(30'h1472b8a5) * $signed(16'h0);
  assign T9179 = T9177[6'h2d:6'h2d];
  assign T9180 = $signed(T9181) / $signed(22'h100000);
  assign T9181 = $signed(31'h435ac1f8) * $signed(16'h1);
  assign twiddle4_3_307_real = T9186 + T9182;
  assign T9182 = {T9185, T9183};
  assign T9183 = $signed(T9184) / $signed(22'h100000);
  assign T9184 = $signed(30'h13e39be9) * $signed(16'h0);
  assign T9185 = T9183[6'h2d:6'h2d];
  assign T9186 = $signed(T9187) / $signed(22'h100000);
  assign T9187 = $signed(31'h432b3c76) * $signed(16'h1);
  assign T9188 = T2943[1'h0:1'h0];
  assign T9189 = T2943[1'h1:1'h1];
  assign T9190 = T9219 ? T9205 : T9191;
  assign T9191 = T9204 ? twiddle4_3_309_real : twiddle4_3_308_real;
  assign twiddle4_3_308_real = T9196 + T9192;
  assign T9192 = {T9195, T9193};
  assign T9193 = $signed(T9194) / $signed(22'h100000);
  assign T9194 = $signed(30'h135410c2) * $signed(16'h0);
  assign T9195 = T9193[6'h2d:6'h2d];
  assign T9196 = $signed(T9197) / $signed(22'h100000);
  assign T9197 = $signed(31'h42fd08aa) * $signed(16'h1);
  assign twiddle4_3_309_real = T9202 + T9198;
  assign T9198 = {T9201, T9199};
  assign T9199 = $signed(T9200) / $signed(22'h100000);
  assign T9200 = $signed(30'h12c41a4e) * $signed(16'h0);
  assign T9201 = T9199[6'h2d:6'h2d];
  assign T9202 = $signed(T9203) / $signed(22'h100000);
  assign T9203 = $signed(31'h42d02794) * $signed(16'h1);
  assign T9204 = T2943[1'h0:1'h0];
  assign T9205 = T9218 ? twiddle4_3_311_real : twiddle4_3_310_real;
  assign twiddle4_3_310_real = T9210 + T9206;
  assign T9206 = {T9209, T9207};
  assign T9207 = $signed(T9208) / $signed(22'h100000);
  assign T9208 = $signed(30'h1233bbab) * $signed(16'h0);
  assign T9209 = T9207[6'h2d:6'h2d];
  assign T9210 = $signed(T9211) / $signed(22'h100000);
  assign T9211 = $signed(31'h42a49a2f) * $signed(16'h1);
  assign twiddle4_3_311_real = T9216 + T9212;
  assign T9212 = {T9215, T9213};
  assign T9213 = $signed(T9214) / $signed(22'h100000);
  assign T9214 = $signed(30'h11a2f7fb) * $signed(16'h0);
  assign T9215 = T9213[6'h2d:6'h2d];
  assign T9216 = $signed(T9217) / $signed(22'h100000);
  assign T9217 = $signed(31'h427a616a) * $signed(16'h1);
  assign T9218 = T2943[1'h0:1'h0];
  assign T9219 = T2943[1'h1:1'h1];
  assign T9220 = T2943[2'h2:2'h2];
  assign T9221 = T9288 ? T9254 : T9222;
  assign T9222 = T9253 ? T9237 : T9223;
  assign T9223 = T9236 ? twiddle4_3_313_real : twiddle4_3_312_real;
  assign twiddle4_3_312_real = T9228 + T9224;
  assign T9224 = {T9227, T9225};
  assign T9225 = $signed(T9226) / $signed(22'h100000);
  assign T9226 = $signed(30'h1111d262) * $signed(16'h0);
  assign T9227 = T9225[6'h2d:6'h2d];
  assign T9228 = $signed(T9229) / $signed(22'h100000);
  assign T9229 = $signed(31'h42517e32) * $signed(16'h1);
  assign twiddle4_3_313_real = T9234 + T9230;
  assign T9230 = {T9233, T9231};
  assign T9231 = $signed(T9232) / $signed(22'h100000);
  assign T9232 = $signed(30'h10804e05) * $signed(16'h0);
  assign T9233 = T9231[6'h2d:6'h2d];
  assign T9234 = $signed(T9235) / $signed(22'h100000);
  assign T9235 = $signed(31'h4229f168) * $signed(16'h1);
  assign T9236 = T2943[1'h0:1'h0];
  assign T9237 = T9252 ? twiddle4_3_315_real : twiddle4_3_314_real;
  assign twiddle4_3_314_real = T9243 + T9238;
  assign T9238 = {T9241, T9239};
  assign T9239 = $signed(T9240) / $signed(22'h100000);
  assign T9240 = $signed(29'hfee6e0d) * $signed(16'h0);
  assign T9241 = T9242 ? 2'h3 : 2'h0;
  assign T9242 = T9239[6'h2c:6'h2c];
  assign T9243 = $signed(T9244) / $signed(22'h100000);
  assign T9244 = $signed(31'h4203bbe8) * $signed(16'h1);
  assign twiddle4_3_315_real = T9250 + T9245;
  assign T9245 = {T9248, T9246};
  assign T9246 = $signed(T9247) / $signed(22'h100000);
  assign T9247 = $signed(29'hf5c35a3) * $signed(16'h0);
  assign T9248 = T9249 ? 2'h3 : 2'h0;
  assign T9249 = T9246[6'h2c:6'h2c];
  assign T9250 = $signed(T9251) / $signed(22'h100000);
  assign T9251 = $signed(31'h41dede87) * $signed(16'h1);
  assign T9252 = T2943[1'h0:1'h0];
  assign T9253 = T2943[1'h1:1'h1];
  assign T9254 = T9287 ? T9271 : T9255;
  assign T9255 = T9270 ? twiddle4_3_317_real : twiddle4_3_316_real;
  assign twiddle4_3_316_real = T9261 + T9256;
  assign T9256 = {T9259, T9257};
  assign T9257 = $signed(T9258) / $signed(22'h100000);
  assign T9258 = $signed(29'hec9a7f2) * $signed(16'h0);
  assign T9259 = T9260 ? 2'h3 : 2'h0;
  assign T9260 = T9257[6'h2c:6'h2c];
  assign T9261 = $signed(T9262) / $signed(22'h100000);
  assign T9262 = $signed(31'h41bb5a12) * $signed(16'h1);
  assign twiddle4_3_317_real = T9268 + T9263;
  assign T9263 = {T9266, T9264};
  assign T9264 = $signed(T9265) / $signed(22'h100000);
  assign T9265 = $signed(29'he36c829) * $signed(16'h0);
  assign T9266 = T9267 ? 2'h3 : 2'h0;
  assign T9267 = T9264[6'h2c:6'h2c];
  assign T9268 = $signed(T9269) / $signed(22'h100000);
  assign T9269 = $signed(31'h41992f4c) * $signed(16'h1);
  assign T9270 = T2943[1'h0:1'h0];
  assign T9271 = T9286 ? twiddle4_3_319_real : twiddle4_3_318_real;
  assign twiddle4_3_318_real = T9277 + T9272;
  assign T9272 = {T9275, T9273};
  assign T9273 = $signed(T9274) / $signed(22'h100000);
  assign T9274 = $signed(29'hda39977) * $signed(16'h0);
  assign T9275 = T9276 ? 2'h3 : 2'h0;
  assign T9276 = T9273[6'h2c:6'h2c];
  assign T9277 = $signed(T9278) / $signed(22'h100000);
  assign T9278 = $signed(31'h41785ef5) * $signed(16'h1);
  assign twiddle4_3_319_real = T9284 + T9279;
  assign T9279 = {T9282, T9280};
  assign T9280 = $signed(T9281) / $signed(22'h100000);
  assign T9281 = $signed(29'hd101f0d) * $signed(16'h0);
  assign T9282 = T9283 ? 2'h3 : 2'h0;
  assign T9283 = T9280[6'h2c:6'h2c];
  assign T9284 = $signed(T9285) / $signed(22'h100000);
  assign T9285 = $signed(31'h4158e9c1) * $signed(16'h1);
  assign T9286 = T2943[1'h0:1'h0];
  assign T9287 = T2943[1'h1:1'h1];
  assign T9288 = T2943[2'h2:2'h2];
  assign T9289 = T2943[2'h3:2'h3];
  assign T9290 = T2943[3'h4:3'h4];
  assign T9291 = T2943[3'h5:3'h5];
  assign T9292 = T9850 ? T9579 : T9293;
  assign T9293 = T9578 ? T9436 : T9294;
  assign T9294 = T9435 ? T9365 : T9295;
  assign T9295 = T9364 ? T9330 : T9296;
  assign T9296 = T9329 ? T9313 : T9297;
  assign T9297 = T9312 ? twiddle4_3_321_real : twiddle4_3_320_real;
  assign twiddle4_3_320_real = T9303 + T9298;
  assign T9298 = {T9301, T9299};
  assign T9299 = $signed(T9300) / $signed(22'h100000);
  assign T9300 = $signed(29'hc7c5c1e) * $signed(16'h0);
  assign T9301 = T9302 ? 2'h3 : 2'h0;
  assign T9302 = T9299[6'h2c:6'h2c];
  assign T9303 = $signed(T9304) / $signed(22'h100000);
  assign T9304 = $signed(31'h413ad061) * $signed(16'h1);
  assign twiddle4_3_321_real = T9310 + T9305;
  assign T9305 = {T9308, T9306};
  assign T9306 = $signed(T9307) / $signed(22'h100000);
  assign T9307 = $signed(29'hbe853dd) * $signed(16'h0);
  assign T9308 = T9309 ? 2'h3 : 2'h0;
  assign T9309 = T9306[6'h2c:6'h2c];
  assign T9310 = $signed(T9311) / $signed(22'h100000);
  assign T9311 = $signed(31'h411e137a) * $signed(16'h1);
  assign T9312 = T2943[1'h0:1'h0];
  assign T9313 = T9328 ? twiddle4_3_323_real : twiddle4_3_322_real;
  assign twiddle4_3_322_real = T9319 + T9314;
  assign T9314 = {T9317, T9315};
  assign T9315 = $signed(T9316) / $signed(22'h100000);
  assign T9316 = $signed(29'hb540982) * $signed(16'h0);
  assign T9317 = T9318 ? 2'h3 : 2'h0;
  assign T9318 = T9315[6'h2c:6'h2c];
  assign T9319 = $signed(T9320) / $signed(22'h100000);
  assign T9320 = $signed(31'h4102b3ad) * $signed(16'h1);
  assign twiddle4_3_323_real = T9326 + T9321;
  assign T9321 = {T9324, T9322};
  assign T9322 = $signed(T9323) / $signed(22'h100000);
  assign T9323 = $signed(29'habf8043) * $signed(16'h0);
  assign T9324 = T9325 ? 2'h3 : 2'h0;
  assign T9325 = T9322[6'h2c:6'h2c];
  assign T9326 = $signed(T9327) / $signed(22'h100000);
  assign T9327 = $signed(31'h40e8b191) * $signed(16'h1);
  assign T9328 = T2943[1'h0:1'h0];
  assign T9329 = T2943[1'h1:1'h1];
  assign T9330 = T9363 ? T9347 : T9331;
  assign T9331 = T9346 ? twiddle4_3_325_real : twiddle4_3_324_real;
  assign twiddle4_3_324_real = T9337 + T9332;
  assign T9332 = {T9335, T9333};
  assign T9333 = $signed(T9334) / $signed(22'h100000);
  assign T9334 = $signed(29'ha2abb58) * $signed(16'h0);
  assign T9335 = T9336 ? 2'h3 : 2'h0;
  assign T9336 = T9333[6'h2c:6'h2c];
  assign T9337 = $signed(T9338) / $signed(22'h100000);
  assign T9338 = $signed(31'h40d00db7) * $signed(16'h1);
  assign twiddle4_3_325_real = T9344 + T9339;
  assign T9339 = {T9342, T9340};
  assign T9340 = $signed(T9341) / $signed(22'h100000);
  assign T9341 = $signed(29'h995bdfc) * $signed(16'h0);
  assign T9342 = T9343 ? 2'h3 : 2'h0;
  assign T9343 = T9340[6'h2c:6'h2c];
  assign T9344 = $signed(T9345) / $signed(22'h100000);
  assign T9345 = $signed(31'h40b8c8a8) * $signed(16'h1);
  assign T9346 = T2943[1'h0:1'h0];
  assign T9347 = T9362 ? twiddle4_3_327_real : twiddle4_3_326_real;
  assign twiddle4_3_326_real = T9353 + T9348;
  assign T9348 = {T9351, T9349};
  assign T9349 = $signed(T9350) / $signed(22'h100000);
  assign T9350 = $signed(29'h9008b6a) * $signed(16'h0);
  assign T9351 = T9352 ? 2'h3 : 2'h0;
  assign T9352 = T9349[6'h2c:6'h2c];
  assign T9353 = $signed(T9354) / $signed(22'h100000);
  assign T9354 = $signed(31'h40a2e2e4) * $signed(16'h1);
  assign twiddle4_3_327_real = T9360 + T9355;
  assign T9355 = {T9358, T9356};
  assign T9356 = $signed(T9357) / $signed(22'h100000);
  assign T9357 = $signed(29'h86b26de) * $signed(16'h0);
  assign T9358 = T9359 ? 2'h3 : 2'h0;
  assign T9359 = T9356[6'h2c:6'h2c];
  assign T9360 = $signed(T9361) / $signed(22'h100000);
  assign T9361 = $signed(31'h408e5ce6) * $signed(16'h1);
  assign T9362 = T2943[1'h0:1'h0];
  assign T9363 = T2943[1'h1:1'h1];
  assign T9364 = T2943[2'h2:2'h2];
  assign T9365 = T9434 ? T9400 : T9366;
  assign T9366 = T9399 ? T9383 : T9367;
  assign T9367 = T9382 ? twiddle4_3_329_real : twiddle4_3_328_real;
  assign twiddle4_3_328_real = T9373 + T9368;
  assign T9368 = {T9371, T9369};
  assign T9369 = $signed(T9370) / $signed(22'h100000);
  assign T9370 = $signed(28'h7d59395) * $signed(16'h0);
  assign T9371 = T9372 ? 3'h7 : 3'h0;
  assign T9372 = T9369[6'h2b:6'h2b];
  assign T9373 = $signed(T9374) / $signed(22'h100000);
  assign T9374 = $signed(31'h407b371f) * $signed(16'h1);
  assign twiddle4_3_329_real = T9380 + T9375;
  assign T9375 = {T9378, T9376};
  assign T9376 = $signed(T9377) / $signed(22'h100000);
  assign T9377 = $signed(28'h73fd4ce) * $signed(16'h0);
  assign T9378 = T9379 ? 3'h7 : 3'h0;
  assign T9379 = T9376[6'h2b:6'h2b];
  assign T9380 = $signed(T9381) / $signed(22'h100000);
  assign T9381 = $signed(31'h406971f9) * $signed(16'h1);
  assign T9382 = T2943[1'h0:1'h0];
  assign T9383 = T9398 ? twiddle4_3_331_real : twiddle4_3_330_real;
  assign twiddle4_3_330_real = T9389 + T9384;
  assign T9384 = {T9387, T9385};
  assign T9385 = $signed(T9386) / $signed(22'h100000);
  assign T9386 = $signed(28'h6a9edc9) * $signed(16'h0);
  assign T9387 = T9388 ? 3'h7 : 3'h0;
  assign T9388 = T9385[6'h2b:6'h2b];
  assign T9389 = $signed(T9390) / $signed(22'h100000);
  assign T9390 = $signed(31'h40590dd8) * $signed(16'h1);
  assign twiddle4_3_331_real = T9396 + T9391;
  assign T9391 = {T9394, T9392};
  assign T9392 = $signed(T9393) / $signed(22'h100000);
  assign T9393 = $signed(28'h613e1c4) * $signed(16'h0);
  assign T9394 = T9395 ? 3'h7 : 3'h0;
  assign T9395 = T9392[6'h2b:6'h2b];
  assign T9396 = $signed(T9397) / $signed(22'h100000);
  assign T9397 = $signed(31'h404a0b16) * $signed(16'h1);
  assign T9398 = T2943[1'h0:1'h0];
  assign T9399 = T2943[1'h1:1'h1];
  assign T9400 = T9433 ? T9417 : T9401;
  assign T9401 = T9416 ? twiddle4_3_333_real : twiddle4_3_332_real;
  assign twiddle4_3_332_real = T9407 + T9402;
  assign T9402 = {T9405, T9403};
  assign T9403 = $signed(T9404) / $signed(22'h100000);
  assign T9404 = $signed(28'h57db402) * $signed(16'h0);
  assign T9405 = T9406 ? 3'h7 : 3'h0;
  assign T9406 = T9403[6'h2b:6'h2b];
  assign T9407 = $signed(T9408) / $signed(22'h100000);
  assign T9408 = $signed(31'h403c6a07) * $signed(16'h1);
  assign twiddle4_3_333_real = T9414 + T9409;
  assign T9409 = {T9412, T9410};
  assign T9410 = $signed(T9411) / $signed(22'h100000);
  assign T9411 = $signed(28'h4e767c4) * $signed(16'h0);
  assign T9412 = T9413 ? 3'h7 : 3'h0;
  assign T9413 = T9410[6'h2b:6'h2b];
  assign T9414 = $signed(T9415) / $signed(22'h100000);
  assign T9415 = $signed(31'h40302af6) * $signed(16'h1);
  assign T9416 = T2943[1'h0:1'h0];
  assign T9417 = T9432 ? twiddle4_3_335_real : twiddle4_3_334_real;
  assign twiddle4_3_334_real = T9423 + T9418;
  assign T9418 = {T9421, T9419};
  assign T9419 = $signed(T9420) / $signed(22'h100000);
  assign T9420 = $signed(28'h451004d) * $signed(16'h0);
  assign T9421 = T9422 ? 3'h7 : 3'h0;
  assign T9422 = T9419[6'h2b:6'h2b];
  assign T9423 = $signed(T9424) / $signed(22'h100000);
  assign T9424 = $signed(31'h40254e27) * $signed(16'h1);
  assign twiddle4_3_335_real = T9430 + T9425;
  assign T9425 = {T9428, T9426};
  assign T9426 = $signed(T9427) / $signed(22'h100000);
  assign T9427 = $signed(27'h3ba80df) * $signed(16'h0);
  assign T9428 = T9429 ? 4'hf : 4'h0;
  assign T9429 = T9426[6'h2a:6'h2a];
  assign T9430 = $signed(T9431) / $signed(22'h100000);
  assign T9431 = $signed(31'h401bd3d7) * $signed(16'h1);
  assign T9432 = T2943[1'h0:1'h0];
  assign T9433 = T2943[1'h1:1'h1];
  assign T9434 = T2943[2'h2:2'h2];
  assign T9435 = T2943[2'h3:2'h3];
  assign T9436 = T9577 ? T9507 : T9437;
  assign T9437 = T9506 ? T9472 : T9438;
  assign T9438 = T9471 ? T9455 : T9439;
  assign T9439 = T9454 ? twiddle4_3_337_real : twiddle4_3_336_real;
  assign twiddle4_3_336_real = T9445 + T9440;
  assign T9440 = {T9443, T9441};
  assign T9441 = $signed(T9442) / $signed(22'h100000);
  assign T9442 = $signed(27'h323ecbe) * $signed(16'h0);
  assign T9443 = T9444 ? 4'hf : 4'h0;
  assign T9444 = T9441[6'h2a:6'h2a];
  assign T9445 = $signed(T9446) / $signed(22'h100000);
  assign T9446 = $signed(31'h4013bc3a) * $signed(16'h1);
  assign twiddle4_3_337_real = T9452 + T9447;
  assign T9447 = {T9450, T9448};
  assign T9448 = $signed(T9449) / $signed(22'h100000);
  assign T9449 = $signed(27'h28d472d) * $signed(16'h0);
  assign T9450 = T9451 ? 4'hf : 4'h0;
  assign T9451 = T9448[6'h2a:6'h2a];
  assign T9452 = $signed(T9453) / $signed(22'h100000);
  assign T9453 = $signed(31'h400d077c) * $signed(16'h1);
  assign T9454 = T2943[1'h0:1'h0];
  assign T9455 = T9470 ? twiddle4_3_339_real : twiddle4_3_338_real;
  assign twiddle4_3_338_real = T9461 + T9456;
  assign T9456 = {T9459, T9457};
  assign T9457 = $signed(T9458) / $signed(22'h100000);
  assign T9458 = $signed(26'h1f69373) * $signed(16'h0);
  assign T9459 = T9460 ? 5'h1f : 5'h0;
  assign T9460 = T9457[6'h29:6'h29];
  assign T9461 = $signed(T9462) / $signed(22'h100000);
  assign T9462 = $signed(31'h4007b5c5) * $signed(16'h1);
  assign twiddle4_3_339_real = T9468 + T9463;
  assign T9463 = {T9466, T9464};
  assign T9464 = $signed(T9465) / $signed(22'h100000);
  assign T9465 = $signed(26'h15fd4d2) * $signed(16'h0);
  assign T9466 = T9467 ? 5'h1f : 5'h0;
  assign T9467 = T9464[6'h29:6'h29];
  assign T9468 = $signed(T9469) / $signed(22'h100000);
  assign T9469 = $signed(31'h4003c730) * $signed(16'h1);
  assign T9470 = T2943[1'h0:1'h0];
  assign T9471 = T2943[1'h1:1'h1];
  assign T9472 = T9505 ? T9489 : T9473;
  assign T9473 = T9488 ? twiddle4_3_341_real : twiddle4_3_340_real;
  assign twiddle4_3_340_real = T9479 + T9474;
  assign T9474 = {T9477, T9475};
  assign T9475 = $signed(T9476) / $signed(22'h100000);
  assign T9476 = $signed(25'hc90e8f) * $signed(16'h0);
  assign T9477 = T9478 ? 6'h3f : 6'h0;
  assign T9478 = T9475[6'h28:6'h28];
  assign T9479 = $signed(T9480) / $signed(22'h100000);
  assign T9480 = $signed(31'h40013bd3) * $signed(16'h1);
  assign twiddle4_3_341_real = T9486 + T9481;
  assign T9481 = {T9484, T9482};
  assign T9482 = $signed(T9483) / $signed(22'h100000);
  assign T9483 = $signed(23'h3243f1) * $signed(16'h0);
  assign T9484 = T9485 ? 8'hff : 8'h0;
  assign T9485 = T9482[6'h26:6'h26];
  assign T9486 = $signed(T9487) / $signed(22'h100000);
  assign T9487 = $signed(31'h400013be) * $signed(16'h1);
  assign T9488 = T2943[1'h0:1'h0];
  assign T9489 = T9504 ? twiddle4_3_343_real : twiddle4_3_342_real;
  assign twiddle4_3_342_real = T9495 + T9490;
  assign T9490 = {T9493, T9491};
  assign T9491 = $signed(T9492) / $signed(22'h100000);
  assign T9492 = $signed(24'h9b783d) * $signed(16'h0);
  assign T9493 = T9494 ? 7'h7f : 7'h0;
  assign T9494 = T9491[6'h27:6'h27];
  assign T9495 = $signed(T9496) / $signed(22'h100000);
  assign T9496 = $signed(31'h40004ef5) * $signed(16'h1);
  assign twiddle4_3_343_real = T9502 + T9497;
  assign T9497 = {T9500, T9498};
  assign T9498 = $signed(T9499) / $signed(22'h100000);
  assign T9499 = $signed(25'h104aeb5) * $signed(16'h0);
  assign T9500 = T9501 ? 6'h3f : 6'h0;
  assign T9501 = T9498[6'h28:6'h28];
  assign T9502 = $signed(T9503) / $signed(22'h100000);
  assign T9503 = $signed(31'h4001ed79) * $signed(16'h1);
  assign T9504 = T2943[1'h0:1'h0];
  assign T9505 = T2943[1'h1:1'h1];
  assign T9506 = T2943[2'h2:2'h2];
  assign T9507 = T9576 ? T9542 : T9508;
  assign T9508 = T9541 ? T9525 : T9509;
  assign T9509 = T9524 ? twiddle4_3_345_real : twiddle4_3_344_real;
  assign twiddle4_3_344_real = T9515 + T9510;
  assign T9510 = {T9513, T9511};
  assign T9511 = $signed(T9512) / $signed(22'h100000);
  assign T9512 = $signed(26'h26deaa1) * $signed(16'h0);
  assign T9513 = T9514 ? 5'h1f : 5'h0;
  assign T9514 = T9511[6'h29:6'h29];
  assign T9515 = $signed(T9516) / $signed(22'h100000);
  assign T9516 = $signed(31'h4004ef3f) * $signed(16'h1);
  assign twiddle4_3_345_real = T9522 + T9517;
  assign T9517 = {T9520, T9518};
  assign T9518 = $signed(T9519) / $signed(22'h100000);
  assign T9519 = $signed(27'h5d72f45) * $signed(16'h0);
  assign T9520 = T9521 ? 4'hf : 4'h0;
  assign T9521 = T9518[6'h2a:6'h2a];
  assign T9522 = $signed(T9523) / $signed(22'h100000);
  assign T9523 = $signed(31'h40095438) * $signed(16'h1);
  assign T9524 = T2943[1'h0:1'h0];
  assign T9525 = T9540 ? twiddle4_3_347_real : twiddle4_3_346_real;
  assign twiddle4_3_346_real = T9531 + T9526;
  assign T9526 = {T9529, T9527};
  assign T9527 = $signed(T9528) / $signed(22'h100000);
  assign T9528 = $signed(27'h5407fe6) * $signed(16'h0);
  assign T9529 = T9530 ? 4'hf : 4'h0;
  assign T9530 = T9527[6'h2a:6'h2a];
  assign T9531 = $signed(T9532) / $signed(22'h100000);
  assign T9532 = $signed(31'h400f1c4b) * $signed(16'h1);
  assign twiddle4_3_347_real = T9538 + T9533;
  assign T9533 = {T9536, T9534};
  assign T9534 = $signed(T9535) / $signed(22'h100000);
  assign T9535 = $signed(27'h4a9dfc9) * $signed(16'h0);
  assign T9536 = T9537 ? 4'hf : 4'h0;
  assign T9537 = T9534[6'h2a:6'h2a];
  assign T9538 = $signed(T9539) / $signed(22'h100000);
  assign T9539 = $signed(31'h40164757) * $signed(16'h1);
  assign T9540 = T2943[1'h0:1'h0];
  assign T9541 = T2943[1'h1:1'h1];
  assign T9542 = T9575 ? T9559 : T9543;
  assign T9543 = T9558 ? twiddle4_3_349_real : twiddle4_3_348_real;
  assign twiddle4_3_348_real = T9549 + T9544;
  assign T9544 = {T9547, T9545};
  assign T9545 = $signed(T9546) / $signed(22'h100000);
  assign T9546 = $signed(27'h4135231) * $signed(16'h0);
  assign T9547 = T9548 ? 4'hf : 4'h0;
  assign T9548 = T9545[6'h2a:6'h2a];
  assign T9549 = $signed(T9550) / $signed(22'h100000);
  assign T9550 = $signed(31'h401ed535) * $signed(16'h1);
  assign twiddle4_3_349_real = T9556 + T9551;
  assign T9551 = {T9554, T9552};
  assign T9552 = $signed(T9553) / $signed(22'h100000);
  assign T9553 = $signed(28'hb7cda63) * $signed(16'h0);
  assign T9554 = T9555 ? 3'h7 : 3'h0;
  assign T9555 = T9552[6'h2b:6'h2b];
  assign T9556 = $signed(T9557) / $signed(22'h100000);
  assign T9557 = $signed(31'h4028c5b6) * $signed(16'h1);
  assign T9558 = T2943[1'h0:1'h0];
  assign T9559 = T9574 ? twiddle4_3_351_real : twiddle4_3_350_real;
  assign twiddle4_3_350_real = T9565 + T9560;
  assign T9560 = {T9563, T9561};
  assign T9561 = $signed(T9562) / $signed(22'h100000);
  assign T9562 = $signed(28'hae67ba2) * $signed(16'h0);
  assign T9563 = T9564 ? 3'h7 : 3'h0;
  assign T9564 = T9561[6'h2b:6'h2b];
  assign T9565 = $signed(T9566) / $signed(22'h100000);
  assign T9566 = $signed(31'h403418a2) * $signed(16'h1);
  assign twiddle4_3_351_real = T9572 + T9567;
  assign T9567 = {T9570, T9568};
  assign T9568 = $signed(T9569) / $signed(22'h100000);
  assign T9569 = $signed(28'ha503931) * $signed(16'h0);
  assign T9570 = T9571 ? 3'h7 : 3'h0;
  assign T9571 = T9568[6'h2b:6'h2b];
  assign T9572 = $signed(T9573) / $signed(22'h100000);
  assign T9573 = $signed(31'h4040cdbb) * $signed(16'h1);
  assign T9574 = T2943[1'h0:1'h0];
  assign T9575 = T2943[1'h1:1'h1];
  assign T9576 = T2943[2'h2:2'h2];
  assign T9577 = T2943[2'h3:2'h3];
  assign T9578 = T2943[3'h4:3'h4];
  assign T9579 = T9849 ? T9722 : T9580;
  assign T9580 = T9721 ? T9651 : T9581;
  assign T9581 = T9650 ? T9616 : T9582;
  assign T9582 = T9615 ? T9599 : T9583;
  assign T9583 = T9598 ? twiddle4_3_353_real : twiddle4_3_352_real;
  assign twiddle4_3_352_real = T9589 + T9584;
  assign T9584 = {T9587, T9585};
  assign T9585 = $signed(T9586) / $signed(22'h100000);
  assign T9586 = $signed(28'h9ba1651) * $signed(16'h0);
  assign T9587 = T9588 ? 3'h7 : 3'h0;
  assign T9588 = T9585[6'h2b:6'h2b];
  assign T9589 = $signed(T9590) / $signed(22'h100000);
  assign T9590 = $signed(31'h404ee4b9) * $signed(16'h1);
  assign twiddle4_3_353_real = T9596 + T9591;
  assign T9591 = {T9594, T9592};
  assign T9592 = $signed(T9593) / $signed(22'h100000);
  assign T9593 = $signed(28'h9241645) * $signed(16'h0);
  assign T9594 = T9595 ? 3'h7 : 3'h0;
  assign T9595 = T9592[6'h2b:6'h2b];
  assign T9596 = $signed(T9597) / $signed(22'h100000);
  assign T9597 = $signed(31'h405e5d4f) * $signed(16'h1);
  assign T9598 = T2943[1'h0:1'h0];
  assign T9599 = T9614 ? twiddle4_3_355_real : twiddle4_3_354_real;
  assign twiddle4_3_354_real = T9605 + T9600;
  assign T9600 = {T9603, T9601};
  assign T9601 = $signed(T9602) / $signed(22'h100000);
  assign T9602 = $signed(28'h88e3c4e) * $signed(16'h0);
  assign T9603 = T9604 ? 3'h7 : 3'h0;
  assign T9604 = T9601[6'h2b:6'h2b];
  assign T9605 = $signed(T9606) / $signed(22'h100000);
  assign T9606 = $signed(31'h406f3727) * $signed(16'h1);
  assign twiddle4_3_355_real = T9612 + T9607;
  assign T9607 = {T9610, T9608};
  assign T9608 = $signed(T9609) / $signed(22'h100000);
  assign T9609 = $signed(29'h17f88baa) * $signed(16'h0);
  assign T9610 = T9611 ? 2'h3 : 2'h0;
  assign T9611 = T9608[6'h2c:6'h2c];
  assign T9612 = $signed(T9613) / $signed(22'h100000);
  assign T9613 = $signed(31'h408171e2) * $signed(16'h1);
  assign T9614 = T2943[1'h0:1'h0];
  assign T9615 = T2943[1'h1:1'h1];
  assign T9616 = T9649 ? T9633 : T9617;
  assign T9617 = T9632 ? twiddle4_3_357_real : twiddle4_3_356_real;
  assign twiddle4_3_356_real = T9623 + T9618;
  assign T9618 = {T9621, T9619};
  assign T9619 = $signed(T9620) / $signed(22'h100000);
  assign T9620 = $signed(29'h17630799) * $signed(16'h0);
  assign T9621 = T9622 ? 2'h3 : 2'h0;
  assign T9622 = T9619[6'h2c:6'h2c];
  assign T9623 = $signed(T9624) / $signed(22'h100000);
  assign T9624 = $signed(31'h40950d1d) * $signed(16'h1);
  assign twiddle4_3_357_real = T9630 + T9625;
  assign T9625 = {T9628, T9626};
  assign T9626 = $signed(T9627) / $signed(22'h100000);
  assign T9627 = $signed(29'h16cdb35a) * $signed(16'h0);
  assign T9628 = T9629 ? 2'h3 : 2'h0;
  assign T9629 = T9626[6'h2c:6'h2c];
  assign T9630 = $signed(T9631) / $signed(22'h100000);
  assign T9631 = $signed(31'h40aa086a) * $signed(16'h1);
  assign T9632 = T2943[1'h0:1'h0];
  assign T9633 = T9648 ? twiddle4_3_359_real : twiddle4_3_358_real;
  assign twiddle4_3_358_real = T9639 + T9634;
  assign T9634 = {T9637, T9635};
  assign T9635 = $signed(T9636) / $signed(22'h100000);
  assign T9636 = $signed(29'h16389228) * $signed(16'h0);
  assign T9637 = T9638 ? 2'h3 : 2'h0;
  assign T9638 = T9635[6'h2c:6'h2c];
  assign T9639 = $signed(T9640) / $signed(22'h100000);
  assign T9640 = $signed(31'h40c06355) * $signed(16'h1);
  assign twiddle4_3_359_real = T9646 + T9641;
  assign T9641 = {T9644, T9642};
  assign T9642 = $signed(T9643) / $signed(22'h100000);
  assign T9643 = $signed(29'h15a3a741) * $signed(16'h0);
  assign T9644 = T9645 ? 2'h3 : 2'h0;
  assign T9645 = T9642[6'h2c:6'h2c];
  assign T9646 = $signed(T9647) / $signed(22'h100000);
  assign T9647 = $signed(31'h40d81d61) * $signed(16'h1);
  assign T9648 = T2943[1'h0:1'h0];
  assign T9649 = T2943[1'h1:1'h1];
  assign T9650 = T2943[2'h2:2'h2];
  assign T9651 = T9720 ? T9686 : T9652;
  assign T9652 = T9685 ? T9669 : T9653;
  assign T9653 = T9668 ? twiddle4_3_361_real : twiddle4_3_360_real;
  assign twiddle4_3_360_real = T9659 + T9654;
  assign T9654 = {T9657, T9655};
  assign T9655 = $signed(T9656) / $signed(22'h100000);
  assign T9656 = $signed(29'h150ef5de) * $signed(16'h0);
  assign T9657 = T9658 ? 2'h3 : 2'h0;
  assign T9658 = T9655[6'h2c:6'h2c];
  assign T9659 = $signed(T9660) / $signed(22'h100000);
  assign T9660 = $signed(31'h40f1360c) * $signed(16'h1);
  assign twiddle4_3_361_real = T9666 + T9661;
  assign T9661 = {T9664, T9662};
  assign T9662 = $signed(T9663) / $signed(22'h100000);
  assign T9663 = $signed(29'h147a813a) * $signed(16'h0);
  assign T9664 = T9665 ? 2'h3 : 2'h0;
  assign T9665 = T9662[6'h2c:6'h2c];
  assign T9666 = $signed(T9667) / $signed(22'h100000);
  assign T9667 = $signed(31'h410bacc8) * $signed(16'h1);
  assign T9668 = T2943[1'h0:1'h0];
  assign T9669 = T9684 ? twiddle4_3_363_real : twiddle4_3_362_real;
  assign twiddle4_3_362_real = T9675 + T9670;
  assign T9670 = {T9673, T9671};
  assign T9671 = $signed(T9672) / $signed(22'h100000);
  assign T9672 = $signed(29'h13e64c8c) * $signed(16'h0);
  assign T9673 = T9674 ? 2'h3 : 2'h0;
  assign T9674 = T9671[6'h2c:6'h2c];
  assign T9675 = $signed(T9676) / $signed(22'h100000);
  assign T9676 = $signed(31'h41278105) * $signed(16'h1);
  assign twiddle4_3_363_real = T9682 + T9677;
  assign T9677 = {T9680, T9678};
  assign T9678 = $signed(T9679) / $signed(22'h100000);
  assign T9679 = $signed(29'h13525b0c) * $signed(16'h0);
  assign T9680 = T9681 ? 2'h3 : 2'h0;
  assign T9681 = T9678[6'h2c:6'h2c];
  assign T9682 = $signed(T9683) / $signed(22'h100000);
  assign T9683 = $signed(31'h4144b226) * $signed(16'h1);
  assign T9684 = T2943[1'h0:1'h0];
  assign T9685 = T2943[1'h1:1'h1];
  assign T9686 = T9719 ? T9703 : T9687;
  assign T9687 = T9702 ? twiddle4_3_365_real : twiddle4_3_364_real;
  assign twiddle4_3_364_real = T9693 + T9688;
  assign T9688 = {T9691, T9689};
  assign T9689 = $signed(T9690) / $signed(22'h100000);
  assign T9690 = $signed(29'h12beafee) * $signed(16'h0);
  assign T9691 = T9692 ? 2'h3 : 2'h0;
  assign T9692 = T9689[6'h2c:6'h2c];
  assign T9693 = $signed(T9694) / $signed(22'h100000);
  assign T9694 = $signed(31'h41633f8a) * $signed(16'h1);
  assign twiddle4_3_365_real = T9700 + T9695;
  assign T9695 = {T9698, T9696};
  assign T9696 = $signed(T9697) / $signed(22'h100000);
  assign T9697 = $signed(29'h122b4e66) * $signed(16'h0);
  assign T9698 = T9699 ? 2'h3 : 2'h0;
  assign T9699 = T9696[6'h2c:6'h2c];
  assign T9700 = $signed(T9701) / $signed(22'h100000);
  assign T9701 = $signed(31'h41832888) * $signed(16'h1);
  assign T9702 = T2943[1'h0:1'h0];
  assign T9703 = T9718 ? twiddle4_3_367_real : twiddle4_3_366_real;
  assign twiddle4_3_366_real = T9709 + T9704;
  assign T9704 = {T9707, T9705};
  assign T9705 = $signed(T9706) / $signed(22'h100000);
  assign T9706 = $signed(29'h119839a7) * $signed(16'h0);
  assign T9707 = T9708 ? 2'h3 : 2'h0;
  assign T9708 = T9705[6'h2c:6'h2c];
  assign T9709 = $signed(T9710) / $signed(22'h100000);
  assign T9710 = $signed(31'h41a46c6e) * $signed(16'h1);
  assign twiddle4_3_367_real = T9716 + T9711;
  assign T9711 = {T9714, T9712};
  assign T9712 = $signed(T9713) / $signed(22'h100000);
  assign T9713 = $signed(29'h110574e1) * $signed(16'h0);
  assign T9714 = T9715 ? 2'h3 : 2'h0;
  assign T9715 = T9712[6'h2c:6'h2c];
  assign T9716 = $signed(T9717) / $signed(22'h100000);
  assign T9717 = $signed(31'h41c70a84) * $signed(16'h1);
  assign T9718 = T2943[1'h0:1'h0];
  assign T9719 = T2943[1'h1:1'h1];
  assign T9720 = T2943[2'h2:2'h2];
  assign T9721 = T2943[2'h3:2'h3];
  assign T9722 = T9848 ? T9786 : T9723;
  assign T9723 = T9785 ? T9755 : T9724;
  assign T9724 = T9754 ? T9740 : T9725;
  assign T9725 = T9739 ? twiddle4_3_369_real : twiddle4_3_368_real;
  assign twiddle4_3_368_real = T9731 + T9726;
  assign T9726 = {T9729, T9727};
  assign T9727 = $signed(T9728) / $signed(22'h100000);
  assign T9728 = $signed(29'h10730343) * $signed(16'h0);
  assign T9729 = T9730 ? 2'h3 : 2'h0;
  assign T9730 = T9727[6'h2c:6'h2c];
  assign T9731 = $signed(T9732) / $signed(22'h100000);
  assign T9732 = $signed(31'h41eb0209) * $signed(16'h1);
  assign twiddle4_3_369_real = T9737 + T9733;
  assign T9733 = {T9736, T9734};
  assign T9734 = $signed(T9735) / $signed(22'h100000);
  assign T9735 = $signed(30'h2fe0e7fa) * $signed(16'h0);
  assign T9736 = T9734[6'h2d:6'h2d];
  assign T9737 = $signed(T9738) / $signed(22'h100000);
  assign T9738 = $signed(31'h42105236) * $signed(16'h1);
  assign T9739 = T2943[1'h0:1'h0];
  assign T9740 = T9753 ? twiddle4_3_371_real : twiddle4_3_370_real;
  assign twiddle4_3_370_real = T9745 + T9741;
  assign T9741 = {T9744, T9742};
  assign T9742 = $signed(T9743) / $signed(22'h100000);
  assign T9743 = $signed(30'h2f4f2631) * $signed(16'h0);
  assign T9744 = T9742[6'h2d:6'h2d];
  assign T9745 = $signed(T9746) / $signed(22'h100000);
  assign T9746 = $signed(31'h4236fa3c) * $signed(16'h1);
  assign twiddle4_3_371_real = T9751 + T9747;
  assign T9747 = {T9750, T9748};
  assign T9748 = $signed(T9749) / $signed(22'h100000);
  assign T9749 = $signed(30'h2ebdc111) * $signed(16'h0);
  assign T9750 = T9748[6'h2d:6'h2d];
  assign T9751 = $signed(T9752) / $signed(22'h100000);
  assign T9752 = $signed(31'h425ef943) * $signed(16'h1);
  assign T9753 = T2943[1'h0:1'h0];
  assign T9754 = T2943[1'h1:1'h1];
  assign T9755 = T9784 ? T9770 : T9756;
  assign T9756 = T9769 ? twiddle4_3_373_real : twiddle4_3_372_real;
  assign twiddle4_3_372_real = T9761 + T9757;
  assign T9757 = {T9760, T9758};
  assign T9758 = $signed(T9759) / $signed(22'h100000);
  assign T9759 = $signed(30'h2e2cbbc1) * $signed(16'h0);
  assign T9760 = T9758[6'h2d:6'h2d];
  assign T9761 = $signed(T9762) / $signed(22'h100000);
  assign T9762 = $signed(31'h42884e6f) * $signed(16'h1);
  assign twiddle4_3_373_real = T9767 + T9763;
  assign T9763 = {T9766, T9764};
  assign T9764 = $signed(T9765) / $signed(22'h100000);
  assign T9765 = $signed(30'h2d9c1967) * $signed(16'h0);
  assign T9766 = T9764[6'h2d:6'h2d];
  assign T9767 = $signed(T9768) / $signed(22'h100000);
  assign T9768 = $signed(31'h42b2f8d9) * $signed(16'h1);
  assign T9769 = T2943[1'h0:1'h0];
  assign T9770 = T9783 ? twiddle4_3_375_real : twiddle4_3_374_real;
  assign twiddle4_3_374_real = T9775 + T9771;
  assign T9771 = {T9774, T9772};
  assign T9772 = $signed(T9773) / $signed(22'h100000);
  assign T9773 = $signed(30'h2d0bdd26) * $signed(16'h0);
  assign T9774 = T9772[6'h2d:6'h2d];
  assign T9775 = $signed(T9776) / $signed(22'h100000);
  assign T9776 = $signed(31'h42def794) * $signed(16'h1);
  assign twiddle4_3_375_real = T9781 + T9777;
  assign T9777 = {T9780, T9778};
  assign T9778 = $signed(T9779) / $signed(22'h100000);
  assign T9779 = $signed(30'h2c7c0a1d) * $signed(16'h0);
  assign T9780 = T9778[6'h2d:6'h2d];
  assign T9781 = $signed(T9782) / $signed(22'h100000);
  assign T9782 = $signed(31'h430c49ad) * $signed(16'h1);
  assign T9783 = T2943[1'h0:1'h0];
  assign T9784 = T2943[1'h1:1'h1];
  assign T9785 = T2943[2'h2:2'h2];
  assign T9786 = T9847 ? T9817 : T9787;
  assign T9787 = T9816 ? T9802 : T9788;
  assign T9788 = T9801 ? twiddle4_3_377_real : twiddle4_3_376_real;
  assign twiddle4_3_376_real = T9793 + T9789;
  assign T9789 = {T9792, T9790};
  assign T9790 = $signed(T9791) / $signed(22'h100000);
  assign T9791 = $signed(30'h2beca36c) * $signed(16'h0);
  assign T9792 = T9790[6'h2d:6'h2d];
  assign T9793 = $signed(T9794) / $signed(22'h100000);
  assign T9794 = $signed(31'h433aee28) * $signed(16'h1);
  assign twiddle4_3_377_real = T9799 + T9795;
  assign T9795 = {T9798, T9796};
  assign T9796 = $signed(T9797) / $signed(22'h100000);
  assign T9797 = $signed(30'h2b5dac2f) * $signed(16'h0);
  assign T9798 = T9796[6'h2d:6'h2d];
  assign T9799 = $signed(T9800) / $signed(22'h100000);
  assign T9800 = $signed(31'h436ae401) * $signed(16'h1);
  assign T9801 = T2943[1'h0:1'h0];
  assign T9802 = T9815 ? twiddle4_3_379_real : twiddle4_3_378_real;
  assign twiddle4_3_378_real = T9807 + T9803;
  assign T9803 = {T9806, T9804};
  assign T9804 = $signed(T9805) / $signed(22'h100000);
  assign T9805 = $signed(30'h2acf2780) * $signed(16'h0);
  assign T9806 = T9804[6'h2d:6'h2d];
  assign T9807 = $signed(T9808) / $signed(22'h100000);
  assign T9808 = $signed(31'h439c2a30) * $signed(16'h1);
  assign twiddle4_3_379_real = T9813 + T9809;
  assign T9809 = {T9812, T9810};
  assign T9810 = $signed(T9811) / $signed(22'h100000);
  assign T9811 = $signed(30'h2a411875) * $signed(16'h0);
  assign T9812 = T9810[6'h2d:6'h2d];
  assign T9813 = $signed(T9814) / $signed(22'h100000);
  assign T9814 = $signed(31'h43cebfa1) * $signed(16'h1);
  assign T9815 = T2943[1'h0:1'h0];
  assign T9816 = T2943[1'h1:1'h1];
  assign T9817 = T9846 ? T9832 : T9818;
  assign T9818 = T9831 ? twiddle4_3_381_real : twiddle4_3_380_real;
  assign twiddle4_3_380_real = T9823 + T9819;
  assign T9819 = {T9822, T9820};
  assign T9820 = $signed(T9821) / $signed(22'h100000);
  assign T9821 = $signed(30'h29b38223) * $signed(16'h0);
  assign T9822 = T9820[6'h2d:6'h2d];
  assign T9823 = $signed(T9824) / $signed(22'h100000);
  assign T9824 = $signed(31'h4402a33c) * $signed(16'h1);
  assign twiddle4_3_381_real = T9829 + T9825;
  assign T9825 = {T9828, T9826};
  assign T9826 = $signed(T9827) / $signed(22'h100000);
  assign T9827 = $signed(30'h2926679d) * $signed(16'h0);
  assign T9828 = T9826[6'h2d:6'h2d];
  assign T9829 = $signed(T9830) / $signed(22'h100000);
  assign T9830 = $signed(31'h4437d3e2) * $signed(16'h1);
  assign T9831 = T2943[1'h0:1'h0];
  assign T9832 = T9845 ? twiddle4_3_383_real : twiddle4_3_382_real;
  assign twiddle4_3_382_real = T9837 + T9833;
  assign T9833 = {T9836, T9834};
  assign T9834 = $signed(T9835) / $signed(22'h100000);
  assign T9835 = $signed(30'h2899cbf1) * $signed(16'h0);
  assign T9836 = T9834[6'h2d:6'h2d];
  assign T9837 = $signed(T9838) / $signed(22'h100000);
  assign T9838 = $signed(31'h446e506a) * $signed(16'h1);
  assign twiddle4_3_383_real = T9843 + T9839;
  assign T9839 = {T9842, T9840};
  assign T9840 = $signed(T9841) / $signed(22'h100000);
  assign T9841 = $signed(30'h280db22d) * $signed(16'h0);
  assign T9842 = T9840[6'h2d:6'h2d];
  assign T9843 = $signed(T9844) / $signed(22'h100000);
  assign T9844 = $signed(31'h44a617a7) * $signed(16'h1);
  assign T9845 = T2943[1'h0:1'h0];
  assign T9846 = T2943[1'h1:1'h1];
  assign T9847 = T2943[2'h2:2'h2];
  assign T9848 = T2943[2'h3:2'h3];
  assign T9849 = T2943[3'h4:3'h4];
  assign T9850 = T2943[3'h5:3'h5];
  assign T9851 = T2943[3'h6:3'h6];
  assign T9852 = T10786 ? T10265 : T9853;
  assign T9853 = T10264 ? T10074 : T9854;
  assign T9854 = T10073 ? T9979 : T9855;
  assign T9855 = T9978 ? T9918 : T9856;
  assign T9856 = T9917 ? T9887 : T9857;
  assign T9857 = T9886 ? T9872 : T9858;
  assign T9858 = T9871 ? twiddle4_3_385_real : twiddle4_3_384_real;
  assign twiddle4_3_384_real = T9863 + T9859;
  assign T9859 = {T9862, T9860};
  assign T9860 = $signed(T9861) / $signed(22'h100000);
  assign T9861 = $signed(30'h27821d5a) * $signed(16'h0);
  assign T9862 = T9860[6'h2d:6'h2d];
  assign T9863 = $signed(T9864) / $signed(22'h100000);
  assign T9864 = $signed(31'h44df2862) * $signed(16'h1);
  assign twiddle4_3_385_real = T9869 + T9865;
  assign T9865 = {T9868, T9866};
  assign T9866 = $signed(T9867) / $signed(22'h100000);
  assign T9867 = $signed(30'h26f7107f) * $signed(16'h0);
  assign T9868 = T9866[6'h2d:6'h2d];
  assign T9869 = $signed(T9870) / $signed(22'h100000);
  assign T9870 = $signed(31'h4519815f) * $signed(16'h1);
  assign T9871 = T2943[1'h0:1'h0];
  assign T9872 = T9885 ? twiddle4_3_387_real : twiddle4_3_386_real;
  assign twiddle4_3_386_real = T9877 + T9873;
  assign T9873 = {T9876, T9874};
  assign T9874 = $signed(T9875) / $signed(22'h100000);
  assign T9875 = $signed(30'h266c8e9f) * $signed(16'h0);
  assign T9876 = T9874[6'h2d:6'h2d];
  assign T9877 = $signed(T9878) / $signed(22'h100000);
  assign T9878 = $signed(31'h4555215b) * $signed(16'h1);
  assign twiddle4_3_387_real = T9883 + T9879;
  assign T9879 = {T9882, T9880};
  assign T9880 = $signed(T9881) / $signed(22'h100000);
  assign T9881 = $signed(30'h25e29abd) * $signed(16'h0);
  assign T9882 = T9880[6'h2d:6'h2d];
  assign T9883 = $signed(T9884) / $signed(22'h100000);
  assign T9884 = $signed(31'h45920709) * $signed(16'h1);
  assign T9885 = T2943[1'h0:1'h0];
  assign T9886 = T2943[1'h1:1'h1];
  assign T9887 = T9916 ? T9902 : T9888;
  assign T9888 = T9901 ? twiddle4_3_389_real : twiddle4_3_388_real;
  assign twiddle4_3_388_real = T9893 + T9889;
  assign T9889 = {T9892, T9890};
  assign T9890 = $signed(T9891) / $signed(22'h100000);
  assign T9891 = $signed(30'h255937d5) * $signed(16'h0);
  assign T9892 = T9890[6'h2d:6'h2d];
  assign T9893 = $signed(T9894) / $signed(22'h100000);
  assign T9894 = $signed(31'h45d03118) * $signed(16'h1);
  assign twiddle4_3_389_real = T9899 + T9895;
  assign T9895 = {T9898, T9896};
  assign T9896 = $signed(T9897) / $signed(22'h100000);
  assign T9897 = $signed(30'h24d068e3) * $signed(16'h0);
  assign T9898 = T9896[6'h2d:6'h2d];
  assign T9899 = $signed(T9900) / $signed(22'h100000);
  assign T9900 = $signed(31'h460f9e2f) * $signed(16'h1);
  assign T9901 = T2943[1'h0:1'h0];
  assign T9902 = T9915 ? twiddle4_3_391_real : twiddle4_3_390_real;
  assign twiddle4_3_390_real = T9907 + T9903;
  assign T9903 = {T9906, T9904};
  assign T9904 = $signed(T9905) / $signed(22'h100000);
  assign T9905 = $signed(30'h244830dd) * $signed(16'h0);
  assign T9906 = T9904[6'h2d:6'h2d];
  assign T9907 = $signed(T9908) / $signed(22'h100000);
  assign T9908 = $signed(31'h46504ced) * $signed(16'h1);
  assign twiddle4_3_391_real = T9913 + T9909;
  assign T9909 = {T9912, T9910};
  assign T9910 = $signed(T9911) / $signed(22'h100000);
  assign T9911 = $signed(30'h23c092b9) * $signed(16'h0);
  assign T9912 = T9910[6'h2d:6'h2d];
  assign T9913 = $signed(T9914) / $signed(22'h100000);
  assign T9914 = $signed(31'h46923bec) * $signed(16'h1);
  assign T9915 = T2943[1'h0:1'h0];
  assign T9916 = T2943[1'h1:1'h1];
  assign T9917 = T2943[2'h2:2'h2];
  assign T9918 = T9977 ? T9949 : T9919;
  assign T9919 = T9948 ? T9934 : T9920;
  assign T9920 = T9933 ? twiddle4_3_393_real : twiddle4_3_392_real;
  assign twiddle4_3_392_real = T9925 + T9921;
  assign T9921 = {T9924, T9922};
  assign T9922 = $signed(T9923) / $signed(22'h100000);
  assign T9923 = $signed(30'h23399167) * $signed(16'h0);
  assign T9924 = T9922[6'h2d:6'h2d];
  assign T9925 = $signed(T9926) / $signed(22'h100000);
  assign T9926 = $signed(31'h46d569be) * $signed(16'h1);
  assign twiddle4_3_393_real = T9931 + T9927;
  assign T9927 = {T9930, T9928};
  assign T9928 = $signed(T9929) / $signed(22'h100000);
  assign T9929 = $signed(30'h22b32fd5) * $signed(16'h0);
  assign T9930 = T9928[6'h2d:6'h2d];
  assign T9931 = $signed(T9932) / $signed(22'h100000);
  assign T9932 = $signed(31'h4719d4ed) * $signed(16'h1);
  assign T9933 = T2943[1'h0:1'h0];
  assign T9934 = T9947 ? twiddle4_3_395_real : twiddle4_3_394_real;
  assign twiddle4_3_394_real = T9939 + T9935;
  assign T9935 = {T9938, T9936};
  assign T9936 = $signed(T9937) / $signed(22'h100000);
  assign T9937 = $signed(30'h222d70ec) * $signed(16'h0);
  assign T9938 = T9936[6'h2d:6'h2d];
  assign T9939 = $signed(T9940) / $signed(22'h100000);
  assign T9940 = $signed(31'h475f7bfe) * $signed(16'h1);
  assign twiddle4_3_395_real = T9945 + T9941;
  assign T9941 = {T9944, T9942};
  assign T9942 = $signed(T9943) / $signed(22'h100000);
  assign T9943 = $signed(30'h21a85793) * $signed(16'h0);
  assign T9944 = T9942[6'h2d:6'h2d];
  assign T9945 = $signed(T9946) / $signed(22'h100000);
  assign T9946 = $signed(31'h47a65d6e) * $signed(16'h1);
  assign T9947 = T2943[1'h0:1'h0];
  assign T9948 = T2943[1'h1:1'h1];
  assign T9949 = T9976 ? T9964 : T9950;
  assign T9950 = T9963 ? twiddle4_3_397_real : twiddle4_3_396_real;
  assign twiddle4_3_396_real = T9955 + T9951;
  assign T9951 = {T9954, T9952};
  assign T9952 = $signed(T9953) / $signed(22'h100000);
  assign T9953 = $signed(30'h2123e6ae) * $signed(16'h0);
  assign T9954 = T9952[6'h2d:6'h2d];
  assign T9955 = $signed(T9956) / $signed(22'h100000);
  assign T9956 = $signed(31'h47ee77b4) * $signed(16'h1);
  assign twiddle4_3_397_real = T9961 + T9957;
  assign T9957 = {T9960, T9958};
  assign T9958 = $signed(T9959) / $signed(22'h100000);
  assign T9959 = $signed(30'h20a0211a) * $signed(16'h0);
  assign T9960 = T9958[6'h2d:6'h2d];
  assign T9961 = $signed(T9962) / $signed(22'h100000);
  assign T9962 = $signed(31'h4837c93e) * $signed(16'h1);
  assign T9963 = T2943[1'h0:1'h0];
  assign T9964 = T9975 ? twiddle4_3_399_real : twiddle4_3_398_real;
  assign twiddle4_3_398_real = T9969 + T9965;
  assign T9965 = {T9968, T9966};
  assign T9966 = $signed(T9967) / $signed(22'h100000);
  assign T9967 = $signed(30'h201d09b5) * $signed(16'h0);
  assign T9968 = T9966[6'h2d:6'h2d];
  assign T9969 = $signed(T9970) / $signed(22'h100000);
  assign T9970 = $signed(31'h48825077) * $signed(16'h1);
  assign twiddle4_3_399_real = T9973 + T9971;
  assign T9971 = $signed(T9972) / $signed(22'h100000);
  assign T9972 = $signed(31'h5f9aa355) * $signed(16'h0);
  assign T9973 = $signed(T9974) / $signed(22'h100000);
  assign T9974 = $signed(31'h48ce0bc1) * $signed(16'h1);
  assign T9975 = T2943[1'h0:1'h0];
  assign T9976 = T2943[1'h1:1'h1];
  assign T9977 = T2943[2'h2:2'h2];
  assign T9978 = T2943[2'h3:2'h3];
  assign T9979 = T10072 ? T10026 : T9980;
  assign T9980 = T10025 ? T10003 : T9981;
  assign T9981 = T10002 ? T9992 : T9982;
  assign T9982 = T9991 ? twiddle4_3_401_real : twiddle4_3_400_real;
  assign twiddle4_3_400_real = T9985 + T9983;
  assign T9983 = $signed(T9984) / $signed(22'h100000);
  assign T9984 = $signed(31'h5f18f0ce) * $signed(16'h0);
  assign T9985 = $signed(T9986) / $signed(22'h100000);
  assign T9986 = $signed(31'h491af976) * $signed(16'h1);
  assign twiddle4_3_401_real = T9989 + T9987;
  assign T9987 = $signed(T9988) / $signed(22'h100000);
  assign T9988 = $signed(31'h5e97f4f1) * $signed(16'h0);
  assign T9989 = $signed(T9990) / $signed(22'h100000);
  assign T9990 = $signed(31'h496917ed) * $signed(16'h1);
  assign T9991 = T2943[1'h0:1'h0];
  assign T9992 = T10001 ? twiddle4_3_403_real : twiddle4_3_402_real;
  assign twiddle4_3_402_real = T9995 + T9993;
  assign T9993 = $signed(T9994) / $signed(22'h100000);
  assign T9994 = $signed(31'h5e17b28a) * $signed(16'h0);
  assign T9995 = $signed(T9996) / $signed(22'h100000);
  assign T9996 = $signed(31'h49b86572) * $signed(16'h1);
  assign twiddle4_3_403_real = T9999 + T9997;
  assign T9997 = $signed(T9998) / $signed(22'h100000);
  assign T9998 = $signed(31'h5d982c61) * $signed(16'h0);
  assign T9999 = $signed(T10000) / $signed(22'h100000);
  assign T10000 = $signed(31'h4a08e04f) * $signed(16'h1);
  assign T10001 = T2943[1'h0:1'h0];
  assign T10002 = T2943[1'h1:1'h1];
  assign T10003 = T10024 ? T10014 : T10004;
  assign T10004 = T10013 ? twiddle4_3_405_real : twiddle4_3_404_real;
  assign twiddle4_3_404_real = T10007 + T10005;
  assign T10005 = $signed(T10006) / $signed(22'h100000);
  assign T10006 = $signed(31'h5d196539) * $signed(16'h0);
  assign T10007 = $signed(T10008) / $signed(22'h100000);
  assign T10008 = $signed(31'h4a5a86c4) * $signed(16'h1);
  assign twiddle4_3_405_real = T10011 + T10009;
  assign T10009 = $signed(T10010) / $signed(22'h100000);
  assign T10010 = $signed(31'h5c9b5fd2) * $signed(16'h0);
  assign T10011 = $signed(T10012) / $signed(22'h100000);
  assign T10012 = $signed(31'h4aad570c) * $signed(16'h1);
  assign T10013 = T2943[1'h0:1'h0];
  assign T10014 = T10023 ? twiddle4_3_407_real : twiddle4_3_406_real;
  assign twiddle4_3_406_real = T10017 + T10015;
  assign T10015 = $signed(T10016) / $signed(22'h100000);
  assign T10016 = $signed(31'h5c1e1ee9) * $signed(16'h0);
  assign T10017 = $signed(T10018) / $signed(22'h100000);
  assign T10018 = $signed(31'h4b014f5b) * $signed(16'h1);
  assign twiddle4_3_407_real = T10021 + T10019;
  assign T10019 = $signed(T10020) / $signed(22'h100000);
  assign T10020 = $signed(31'h5ba1a534) * $signed(16'h0);
  assign T10021 = $signed(T10022) / $signed(22'h100000);
  assign T10022 = $signed(31'h4b566ddf) * $signed(16'h1);
  assign T10023 = T2943[1'h0:1'h0];
  assign T10024 = T2943[1'h1:1'h1];
  assign T10025 = T2943[2'h2:2'h2];
  assign T10026 = T10071 ? T10049 : T10027;
  assign T10027 = T10048 ? T10038 : T10028;
  assign T10028 = T10037 ? twiddle4_3_409_real : twiddle4_3_408_real;
  assign twiddle4_3_408_real = T10031 + T10029;
  assign T10029 = $signed(T10030) / $signed(22'h100000);
  assign T10030 = $signed(31'h5b25f567) * $signed(16'h0);
  assign T10031 = $signed(T10032) / $signed(22'h100000);
  assign T10032 = $signed(31'h4bacb0c0) * $signed(16'h1);
  assign twiddle4_3_409_real = T10035 + T10033;
  assign T10033 = $signed(T10034) / $signed(22'h100000);
  assign T10034 = $signed(31'h5aab1230) * $signed(16'h0);
  assign T10035 = $signed(T10036) / $signed(22'h100000);
  assign T10036 = $signed(31'h4c04161e) * $signed(16'h1);
  assign T10037 = T2943[1'h0:1'h0];
  assign T10038 = T10047 ? twiddle4_3_411_real : twiddle4_3_410_real;
  assign twiddle4_3_410_real = T10041 + T10039;
  assign T10039 = $signed(T10040) / $signed(22'h100000);
  assign T10040 = $signed(31'h5a30fe39) * $signed(16'h0);
  assign T10041 = $signed(T10042) / $signed(22'h100000);
  assign T10042 = $signed(31'h4c5c9c15) * $signed(16'h1);
  assign twiddle4_3_411_real = T10045 + T10043;
  assign T10043 = $signed(T10044) / $signed(22'h100000);
  assign T10044 = $signed(31'h59b7bc28) * $signed(16'h0);
  assign T10045 = $signed(T10046) / $signed(22'h100000);
  assign T10046 = $signed(31'h4cb640b8) * $signed(16'h1);
  assign T10047 = T2943[1'h0:1'h0];
  assign T10048 = T2943[1'h1:1'h1];
  assign T10049 = T10070 ? T10060 : T10050;
  assign T10050 = T10059 ? twiddle4_3_413_real : twiddle4_3_412_real;
  assign twiddle4_3_412_real = T10053 + T10051;
  assign T10051 = $signed(T10052) / $signed(22'h100000);
  assign T10052 = $signed(31'h593f4e9e) * $signed(16'h0);
  assign T10053 = $signed(T10054) / $signed(22'h100000);
  assign T10054 = $signed(31'h4d110217) * $signed(16'h1);
  assign twiddle4_3_413_real = T10057 + T10055;
  assign T10055 = $signed(T10056) / $signed(22'h100000);
  assign T10056 = $signed(31'h58c7b839) * $signed(16'h0);
  assign T10057 = $signed(T10058) / $signed(22'h100000);
  assign T10058 = $signed(31'h4d6cde39) * $signed(16'h1);
  assign T10059 = T2943[1'h0:1'h0];
  assign T10060 = T10069 ? twiddle4_3_415_real : twiddle4_3_414_real;
  assign twiddle4_3_414_real = T10063 + T10061;
  assign T10061 = $signed(T10062) / $signed(22'h100000);
  assign T10062 = $signed(31'h5850fb8f) * $signed(16'h0);
  assign T10063 = $signed(T10064) / $signed(22'h100000);
  assign T10064 = $signed(31'h4dc9d321) * $signed(16'h1);
  assign twiddle4_3_415_real = T10067 + T10065;
  assign T10065 = $signed(T10066) / $signed(22'h100000);
  assign T10066 = $signed(31'h57db1b34) * $signed(16'h0);
  assign T10067 = $signed(T10068) / $signed(22'h100000);
  assign T10068 = $signed(31'h4e27deca) * $signed(16'h1);
  assign T10069 = T2943[1'h0:1'h0];
  assign T10070 = T2943[1'h1:1'h1];
  assign T10071 = T2943[2'h2:2'h2];
  assign T10072 = T2943[2'h3:2'h3];
  assign T10073 = T2943[3'h4:3'h4];
  assign T10074 = T10263 ? T10169 : T10075;
  assign T10075 = T10168 ? T10122 : T10076;
  assign T10076 = T10121 ? T10099 : T10077;
  assign T10077 = T10098 ? T10088 : T10078;
  assign T10078 = T10087 ? twiddle4_3_417_real : twiddle4_3_416_real;
  assign twiddle4_3_416_real = T10081 + T10079;
  assign T10079 = $signed(T10080) / $signed(22'h100000);
  assign T10080 = $signed(31'h576619b6) * $signed(16'h0);
  assign T10081 = $signed(T10082) / $signed(22'h100000);
  assign T10082 = $signed(31'h4e86ff2a) * $signed(16'h1);
  assign twiddle4_3_417_real = T10085 + T10083;
  assign T10083 = $signed(T10084) / $signed(22'h100000);
  assign T10084 = $signed(31'h56f1f9a0) * $signed(16'h0);
  assign T10085 = $signed(T10086) / $signed(22'h100000);
  assign T10086 = $signed(31'h4ee73232) * $signed(16'h1);
  assign T10087 = T2943[1'h0:1'h0];
  assign T10088 = T10097 ? twiddle4_3_419_real : twiddle4_3_418_real;
  assign twiddle4_3_418_real = T10091 + T10089;
  assign T10089 = $signed(T10090) / $signed(22'h100000);
  assign T10090 = $signed(31'h567ebd75) * $signed(16'h0);
  assign T10091 = $signed(T10092) / $signed(22'h100000);
  assign T10092 = $signed(31'h4f4875cb) * $signed(16'h1);
  assign twiddle4_3_419_real = T10095 + T10093;
  assign T10093 = $signed(T10094) / $signed(22'h100000);
  assign T10094 = $signed(31'h560c67b5) * $signed(16'h0);
  assign T10095 = $signed(T10096) / $signed(22'h100000);
  assign T10096 = $signed(31'h4faac7d9) * $signed(16'h1);
  assign T10097 = T2943[1'h0:1'h0];
  assign T10098 = T2943[1'h1:1'h1];
  assign T10099 = T10120 ? T10110 : T10100;
  assign T10100 = T10109 ? twiddle4_3_421_real : twiddle4_3_420_real;
  assign twiddle4_3_420_real = T10103 + T10101;
  assign T10101 = $signed(T10102) / $signed(22'h100000);
  assign T10102 = $signed(31'h559afadb) * $signed(16'h0);
  assign T10103 = $signed(T10104) / $signed(22'h100000);
  assign T10104 = $signed(31'h500e263a) * $signed(16'h1);
  assign twiddle4_3_421_real = T10107 + T10105;
  assign T10105 = $signed(T10106) / $signed(22'h100000);
  assign T10106 = $signed(31'h552a795d) * $signed(16'h0);
  assign T10107 = $signed(T10108) / $signed(22'h100000);
  assign T10108 = $signed(31'h50728ec7) * $signed(16'h1);
  assign T10109 = T2943[1'h0:1'h0];
  assign T10110 = T10119 ? twiddle4_3_423_real : twiddle4_3_422_real;
  assign twiddle4_3_422_real = T10113 + T10111;
  assign T10111 = $signed(T10112) / $signed(22'h100000);
  assign T10112 = $signed(31'h54bae5ac) * $signed(16'h0);
  assign T10113 = $signed(T10114) / $signed(22'h100000);
  assign T10114 = $signed(31'h50d7ff52) * $signed(16'h1);
  assign twiddle4_3_423_real = T10117 + T10115;
  assign T10115 = $signed(T10116) / $signed(22'h100000);
  assign T10116 = $signed(31'h544c4232) * $signed(16'h0);
  assign T10117 = $signed(T10118) / $signed(22'h100000);
  assign T10118 = $signed(31'h513e75a8) * $signed(16'h1);
  assign T10119 = T2943[1'h0:1'h0];
  assign T10120 = T2943[1'h1:1'h1];
  assign T10121 = T2943[2'h2:2'h2];
  assign T10122 = T10167 ? T10145 : T10123;
  assign T10123 = T10144 ? T10134 : T10124;
  assign T10124 = T10133 ? twiddle4_3_425_real : twiddle4_3_424_real;
  assign twiddle4_3_424_real = T10127 + T10125;
  assign T10125 = $signed(T10126) / $signed(22'h100000);
  assign T10126 = $signed(31'h53de9156) * $signed(16'h0);
  assign T10127 = $signed(T10128) / $signed(22'h100000);
  assign T10128 = $signed(31'h51a5ef91) * $signed(16'h1);
  assign twiddle4_3_425_real = T10131 + T10129;
  assign T10129 = $signed(T10130) / $signed(22'h100000);
  assign T10130 = $signed(31'h5371d57a) * $signed(16'h0);
  assign T10131 = $signed(T10132) / $signed(22'h100000);
  assign T10132 = $signed(31'h520e6acd) * $signed(16'h1);
  assign T10133 = T2943[1'h0:1'h0];
  assign T10134 = T10143 ? twiddle4_3_427_real : twiddle4_3_426_real;
  assign twiddle4_3_426_real = T10137 + T10135;
  assign T10135 = $signed(T10136) / $signed(22'h100000);
  assign T10136 = $signed(31'h530610f7) * $signed(16'h0);
  assign T10137 = $signed(T10138) / $signed(22'h100000);
  assign T10138 = $signed(31'h5277e519) * $signed(16'h1);
  assign twiddle4_3_427_real = T10141 + T10139;
  assign T10139 = $signed(T10140) / $signed(22'h100000);
  assign T10140 = $signed(31'h529b4626) * $signed(16'h0);
  assign T10141 = $signed(T10142) / $signed(22'h100000);
  assign T10142 = $signed(31'h52e25c2b) * $signed(16'h1);
  assign T10143 = T2943[1'h0:1'h0];
  assign T10144 = T2943[1'h1:1'h1];
  assign T10145 = T10166 ? T10156 : T10146;
  assign T10146 = T10155 ? twiddle4_3_429_real : twiddle4_3_428_real;
  assign twiddle4_3_428_real = T10149 + T10147;
  assign T10147 = $signed(T10148) / $signed(22'h100000);
  assign T10148 = $signed(31'h52317757) * $signed(16'h0);
  assign T10149 = $signed(T10150) / $signed(22'h100000);
  assign T10150 = $signed(31'h534dcdb5) * $signed(16'h1);
  assign twiddle4_3_429_real = T10153 + T10151;
  assign T10151 = $signed(T10152) / $signed(22'h100000);
  assign T10152 = $signed(31'h51c8a6d4) * $signed(16'h0);
  assign T10153 = $signed(T10154) / $signed(22'h100000);
  assign T10154 = $signed(31'h53ba3761) * $signed(16'h1);
  assign T10155 = T2943[1'h0:1'h0];
  assign T10156 = T10165 ? twiddle4_3_431_real : twiddle4_3_430_real;
  assign twiddle4_3_430_real = T10159 + T10157;
  assign T10157 = $signed(T10158) / $signed(22'h100000);
  assign T10158 = $signed(31'h5160d6e5) * $signed(16'h0);
  assign T10159 = $signed(T10160) / $signed(22'h100000);
  assign T10160 = $signed(31'h542796d5) * $signed(16'h1);
  assign twiddle4_3_431_real = T10163 + T10161;
  assign T10161 = $signed(T10162) / $signed(22'h100000);
  assign T10162 = $signed(31'h50fa09c9) * $signed(16'h0);
  assign T10163 = $signed(T10164) / $signed(22'h100000);
  assign T10164 = $signed(31'h5495e9b4) * $signed(16'h1);
  assign T10165 = T2943[1'h0:1'h0];
  assign T10166 = T2943[1'h1:1'h1];
  assign T10167 = T2943[2'h2:2'h2];
  assign T10168 = T2943[2'h3:2'h3];
  assign T10169 = T10262 ? T10216 : T10170;
  assign T10170 = T10215 ? T10193 : T10171;
  assign T10171 = T10192 ? T10182 : T10172;
  assign T10172 = T10181 ? twiddle4_3_433_real : twiddle4_3_432_real;
  assign twiddle4_3_432_real = T10175 + T10173;
  assign T10173 = $signed(T10174) / $signed(22'h100000);
  assign T10174 = $signed(31'h509441bc) * $signed(16'h0);
  assign T10175 = $signed(T10176) / $signed(22'h100000);
  assign T10176 = $signed(31'h55052d97) * $signed(16'h1);
  assign twiddle4_3_433_real = T10179 + T10177;
  assign T10177 = $signed(T10178) / $signed(22'h100000);
  assign T10178 = $signed(31'h502f80f1) * $signed(16'h0);
  assign T10179 = $signed(T10180) / $signed(22'h100000);
  assign T10180 = $signed(31'h55756016) * $signed(16'h1);
  assign T10181 = T2943[1'h0:1'h0];
  assign T10182 = T10191 ? twiddle4_3_435_real : twiddle4_3_434_real;
  assign twiddle4_3_434_real = T10185 + T10183;
  assign T10183 = $signed(T10184) / $signed(22'h100000);
  assign T10184 = $signed(31'h4fcbc999) * $signed(16'h0);
  assign T10185 = $signed(T10186) / $signed(22'h100000);
  assign T10186 = $signed(31'h55e67ec2) * $signed(16'h1);
  assign twiddle4_3_435_real = T10189 + T10187;
  assign T10187 = $signed(T10188) / $signed(22'h100000);
  assign T10188 = $signed(31'h4f691ddd) * $signed(16'h0);
  assign T10189 = $signed(T10190) / $signed(22'h100000);
  assign T10190 = $signed(31'h56588726) * $signed(16'h1);
  assign T10191 = T2943[1'h0:1'h0];
  assign T10192 = T2943[1'h1:1'h1];
  assign T10193 = T10214 ? T10204 : T10194;
  assign T10194 = T10203 ? twiddle4_3_437_real : twiddle4_3_436_real;
  assign twiddle4_3_436_real = T10197 + T10195;
  assign T10195 = $signed(T10196) / $signed(22'h100000);
  assign T10196 = $signed(31'h4f077fe1) * $signed(16'h0);
  assign T10197 = $signed(T10198) / $signed(22'h100000);
  assign T10198 = $signed(31'h56cb76c9) * $signed(16'h1);
  assign twiddle4_3_437_real = T10201 + T10199;
  assign T10199 = $signed(T10200) / $signed(22'h100000);
  assign T10200 = $signed(31'h4ea6f1c3) * $signed(16'h0);
  assign T10201 = $signed(T10202) / $signed(22'h100000);
  assign T10202 = $signed(31'h573f4b2e) * $signed(16'h1);
  assign T10203 = T2943[1'h0:1'h0];
  assign T10204 = T10213 ? twiddle4_3_439_real : twiddle4_3_438_real;
  assign twiddle4_3_438_real = T10207 + T10205;
  assign T10205 = $signed(T10206) / $signed(22'h100000);
  assign T10206 = $signed(31'h4e47759a) * $signed(16'h0);
  assign T10207 = $signed(T10208) / $signed(22'h100000);
  assign T10208 = $signed(31'h57b401d1) * $signed(16'h1);
  assign twiddle4_3_439_real = T10211 + T10209;
  assign T10209 = $signed(T10210) / $signed(22'h100000);
  assign T10210 = $signed(31'h4de90d7a) * $signed(16'h0);
  assign T10211 = $signed(T10212) / $signed(22'h100000);
  assign T10212 = $signed(31'h5829982b) * $signed(16'h1);
  assign T10213 = T2943[1'h0:1'h0];
  assign T10214 = T2943[1'h1:1'h1];
  assign T10215 = T2943[2'h2:2'h2];
  assign T10216 = T10261 ? T10239 : T10217;
  assign T10217 = T10238 ? T10228 : T10218;
  assign T10218 = T10227 ? twiddle4_3_441_real : twiddle4_3_440_real;
  assign twiddle4_3_440_real = T10221 + T10219;
  assign T10219 = $signed(T10220) / $signed(22'h100000);
  assign T10220 = $signed(31'h4d8bbb6d) * $signed(16'h0);
  assign T10221 = $signed(T10222) / $signed(22'h100000);
  assign T10222 = $signed(31'h58a00bae) * $signed(16'h1);
  assign twiddle4_3_441_real = T10225 + T10223;
  assign T10223 = $signed(T10224) / $signed(22'h100000);
  assign T10224 = $signed(31'h4d2f817b) * $signed(16'h0);
  assign T10225 = $signed(T10226) / $signed(22'h100000);
  assign T10226 = $signed(31'h591759c9) * $signed(16'h1);
  assign T10227 = T2943[1'h0:1'h0];
  assign T10228 = T10237 ? twiddle4_3_443_real : twiddle4_3_442_real;
  assign twiddle4_3_442_real = T10231 + T10229;
  assign T10229 = $signed(T10230) / $signed(22'h100000);
  assign T10230 = $signed(31'h4cd461a3) * $signed(16'h0);
  assign T10231 = $signed(T10232) / $signed(22'h100000);
  assign T10232 = $signed(31'h598f7fe6) * $signed(16'h1);
  assign twiddle4_3_443_real = T10235 + T10233;
  assign T10233 = $signed(T10234) / $signed(22'h100000);
  assign T10234 = $signed(31'h4c7a5ddf) * $signed(16'h0);
  assign T10235 = $signed(T10236) / $signed(22'h100000);
  assign T10236 = $signed(31'h5a087b6a) * $signed(16'h1);
  assign T10237 = T2943[1'h0:1'h0];
  assign T10238 = T2943[1'h1:1'h1];
  assign T10239 = T10260 ? T10250 : T10240;
  assign T10240 = T10249 ? twiddle4_3_445_real : twiddle4_3_444_real;
  assign twiddle4_3_444_real = T10243 + T10241;
  assign T10241 = $signed(T10242) / $signed(22'h100000);
  assign T10242 = $signed(31'h4c217822) * $signed(16'h0);
  assign T10243 = $signed(T10244) / $signed(22'h100000);
  assign T10244 = $signed(31'h5a8249b5) * $signed(16'h1);
  assign twiddle4_3_445_real = T10247 + T10245;
  assign T10245 = $signed(T10246) / $signed(22'h100000);
  assign T10246 = $signed(31'h4bc9b25b) * $signed(16'h0);
  assign T10247 = $signed(T10248) / $signed(22'h100000);
  assign T10248 = $signed(31'h5afce822) * $signed(16'h1);
  assign T10249 = T2943[1'h0:1'h0];
  assign T10250 = T10259 ? twiddle4_3_447_real : twiddle4_3_446_real;
  assign twiddle4_3_446_real = T10253 + T10251;
  assign T10251 = $signed(T10252) / $signed(22'h100000);
  assign T10252 = $signed(31'h4b730e70) * $signed(16'h0);
  assign T10253 = $signed(T10254) / $signed(22'h100000);
  assign T10254 = $signed(31'h5b785409) * $signed(16'h1);
  assign twiddle4_3_447_real = T10257 + T10255;
  assign T10255 = $signed(T10256) / $signed(22'h100000);
  assign T10256 = $signed(31'h4b1d8e43) * $signed(16'h0);
  assign T10257 = $signed(T10258) / $signed(22'h100000);
  assign T10258 = $signed(31'h5bf48abe) * $signed(16'h1);
  assign T10259 = T2943[1'h0:1'h0];
  assign T10260 = T2943[1'h1:1'h1];
  assign T10261 = T2943[2'h2:2'h2];
  assign T10262 = T2943[2'h3:2'h3];
  assign T10263 = T2943[3'h4:3'h4];
  assign T10264 = T2943[3'h5:3'h5];
  assign T10265 = T10785 ? T10504 : T10266;
  assign T10266 = T10503 ? T10377 : T10267;
  assign T10267 = T10376 ? T10314 : T10268;
  assign T10268 = T10313 ? T10291 : T10269;
  assign T10269 = T10290 ? T10280 : T10270;
  assign T10270 = T10279 ? twiddle4_3_449_real : twiddle4_3_448_real;
  assign twiddle4_3_448_real = T10273 + T10271;
  assign T10271 = $signed(T10272) / $signed(22'h100000);
  assign T10272 = $signed(31'h4ac933ae) * $signed(16'h0);
  assign T10273 = $signed(T10274) / $signed(22'h100000);
  assign T10274 = $signed(31'h5c71898d) * $signed(16'h1);
  assign twiddle4_3_449_real = T10277 + T10275;
  assign T10275 = $signed(T10276) / $signed(22'h100000);
  assign T10276 = $signed(31'h4a760086) * $signed(16'h0);
  assign T10277 = $signed(T10278) / $signed(22'h100000);
  assign T10278 = $signed(31'h5cef4dc2) * $signed(16'h1);
  assign T10279 = T2943[1'h0:1'h0];
  assign T10280 = T10289 ? twiddle4_3_451_real : twiddle4_3_450_real;
  assign twiddle4_3_450_real = T10283 + T10281;
  assign T10281 = $signed(T10282) / $signed(22'h100000);
  assign T10282 = $signed(31'h4a23f698) * $signed(16'h0);
  assign T10283 = $signed(T10284) / $signed(22'h100000);
  assign T10284 = $signed(31'h5d6dd4a2) * $signed(16'h1);
  assign twiddle4_3_451_real = T10287 + T10285;
  assign T10285 = $signed(T10286) / $signed(22'h100000);
  assign T10286 = $signed(31'h49d317ac) * $signed(16'h0);
  assign T10287 = $signed(T10288) / $signed(22'h100000);
  assign T10288 = $signed(31'h5ded1b6f) * $signed(16'h1);
  assign T10289 = T2943[1'h0:1'h0];
  assign T10290 = T2943[1'h1:1'h1];
  assign T10291 = T10312 ? T10302 : T10292;
  assign T10292 = T10301 ? twiddle4_3_453_real : twiddle4_3_452_real;
  assign twiddle4_3_452_real = T10295 + T10293;
  assign T10293 = $signed(T10294) / $signed(22'h100000);
  assign T10294 = $signed(31'h49836583) * $signed(16'h0);
  assign T10295 = $signed(T10296) / $signed(22'h100000);
  assign T10296 = $signed(31'h5e6d1f66) * $signed(16'h1);
  assign twiddle4_3_453_real = T10299 + T10297;
  assign T10297 = $signed(T10298) / $signed(22'h100000);
  assign T10298 = $signed(31'h4934e1d7) * $signed(16'h0);
  assign T10299 = $signed(T10300) / $signed(22'h100000);
  assign T10300 = $signed(31'h5eedddc0) * $signed(16'h1);
  assign T10301 = T2943[1'h0:1'h0];
  assign T10302 = T10311 ? twiddle4_3_455_real : twiddle4_3_454_real;
  assign twiddle4_3_454_real = T10305 + T10303;
  assign T10303 = $signed(T10304) / $signed(22'h100000);
  assign T10304 = $signed(31'h48e78e5c) * $signed(16'h0);
  assign T10305 = $signed(T10306) / $signed(22'h100000);
  assign T10306 = $signed(31'h5f6f53b3) * $signed(16'h1);
  assign twiddle4_3_455_real = T10309 + T10307;
  assign T10307 = $signed(T10308) / $signed(22'h100000);
  assign T10308 = $signed(31'h489b6cbf) * $signed(16'h0);
  assign T10309 = $signed(T10310) / $signed(22'h100000);
  assign T10310 = $signed(31'h5ff17e70) * $signed(16'h1);
  assign T10311 = T2943[1'h0:1'h0];
  assign T10312 = T2943[1'h1:1'h1];
  assign T10313 = T2943[2'h2:2'h2];
  assign T10314 = T10375 ? T10345 : T10315;
  assign T10315 = T10344 ? T10330 : T10316;
  assign T10316 = T10329 ? twiddle4_3_457_real : twiddle4_3_456_real;
  assign twiddle4_3_456_real = T10319 + T10317;
  assign T10317 = $signed(T10318) / $signed(22'h100000);
  assign T10318 = $signed(31'h48507ea8) * $signed(16'h0);
  assign T10319 = {T10322, T10320};
  assign T10320 = $signed(T10321) / $signed(22'h100000);
  assign T10321 = $signed(30'h20745b25) * $signed(16'h1);
  assign T10322 = T10320[6'h2d:6'h2d];
  assign twiddle4_3_457_real = T10325 + T10323;
  assign T10323 = $signed(T10324) / $signed(22'h100000);
  assign T10324 = $signed(31'h4806c5b5) * $signed(16'h0);
  assign T10325 = {T10328, T10326};
  assign T10326 = $signed(T10327) / $signed(22'h100000);
  assign T10327 = $signed(30'h20f7e6fa) * $signed(16'h1);
  assign T10328 = T10326[6'h2d:6'h2d];
  assign T10329 = T2943[1'h0:1'h0];
  assign T10330 = T10343 ? twiddle4_3_459_real : twiddle4_3_458_real;
  assign twiddle4_3_458_real = T10333 + T10331;
  assign T10331 = $signed(T10332) / $signed(22'h100000);
  assign T10332 = $signed(31'h47be4381) * $signed(16'h0);
  assign T10333 = {T10336, T10334};
  assign T10334 = $signed(T10335) / $signed(22'h100000);
  assign T10335 = $signed(30'h217c1f16) * $signed(16'h1);
  assign T10336 = T10334[6'h2d:6'h2d];
  assign twiddle4_3_459_real = T10339 + T10337;
  assign T10337 = $signed(T10338) / $signed(22'h100000);
  assign T10338 = $signed(31'h4776f99e) * $signed(16'h0);
  assign T10339 = {T10342, T10340};
  assign T10340 = $signed(T10341) / $signed(22'h100000);
  assign T10341 = $signed(30'h2201009a) * $signed(16'h1);
  assign T10342 = T10340[6'h2d:6'h2d];
  assign T10343 = T2943[1'h0:1'h0];
  assign T10344 = T2943[1'h1:1'h1];
  assign T10345 = T10374 ? T10360 : T10346;
  assign T10346 = T10359 ? twiddle4_3_461_real : twiddle4_3_460_real;
  assign twiddle4_3_460_real = T10349 + T10347;
  assign T10347 = $signed(T10348) / $signed(22'h100000);
  assign T10348 = $signed(31'h4730e997) * $signed(16'h0);
  assign T10349 = {T10352, T10350};
  assign T10350 = $signed(T10351) / $signed(22'h100000);
  assign T10351 = $signed(30'h228688a5) * $signed(16'h1);
  assign T10352 = T10350[6'h2d:6'h2d];
  assign twiddle4_3_461_real = T10355 + T10353;
  assign T10353 = $signed(T10354) / $signed(22'h100000);
  assign T10354 = $signed(31'h46ec14f2) * $signed(16'h0);
  assign T10355 = {T10358, T10356};
  assign T10356 = $signed(T10357) / $signed(22'h100000);
  assign T10357 = $signed(30'h230cb452) * $signed(16'h1);
  assign T10358 = T10356[6'h2d:6'h2d];
  assign T10359 = T2943[1'h0:1'h0];
  assign T10360 = T10373 ? twiddle4_3_463_real : twiddle4_3_462_real;
  assign twiddle4_3_462_real = T10363 + T10361;
  assign T10361 = $signed(T10362) / $signed(22'h100000);
  assign T10362 = $signed(31'h46a87d2d) * $signed(16'h0);
  assign T10363 = {T10366, T10364};
  assign T10364 = $signed(T10365) / $signed(22'h100000);
  assign T10365 = $signed(30'h239380b7) * $signed(16'h1);
  assign T10366 = T10364[6'h2d:6'h2d];
  assign twiddle4_3_463_real = T10369 + T10367;
  assign T10367 = $signed(T10368) / $signed(22'h100000);
  assign T10368 = $signed(31'h466623bf) * $signed(16'h0);
  assign T10369 = {T10372, T10370};
  assign T10370 = $signed(T10371) / $signed(22'h100000);
  assign T10371 = $signed(30'h241aeae9) * $signed(16'h1);
  assign T10372 = T10370[6'h2d:6'h2d];
  assign T10373 = T2943[1'h0:1'h0];
  assign T10374 = T2943[1'h1:1'h1];
  assign T10375 = T2943[2'h2:2'h2];
  assign T10376 = T2943[2'h3:2'h3];
  assign T10377 = T10502 ? T10440 : T10378;
  assign T10378 = T10439 ? T10409 : T10379;
  assign T10379 = T10408 ? T10394 : T10380;
  assign T10380 = T10393 ? twiddle4_3_465_real : twiddle4_3_464_real;
  assign twiddle4_3_464_real = T10383 + T10381;
  assign T10381 = $signed(T10382) / $signed(22'h100000);
  assign T10382 = $signed(31'h46250a18) * $signed(16'h0);
  assign T10383 = {T10386, T10384};
  assign T10384 = $signed(T10385) / $signed(22'h100000);
  assign T10385 = $signed(30'h24a2eff7) * $signed(16'h1);
  assign T10386 = T10384[6'h2d:6'h2d];
  assign twiddle4_3_465_real = T10389 + T10387;
  assign T10387 = $signed(T10388) / $signed(22'h100000);
  assign T10388 = $signed(31'h45e531a2) * $signed(16'h0);
  assign T10389 = {T10392, T10390};
  assign T10390 = $signed(T10391) / $signed(22'h100000);
  assign T10391 = $signed(30'h252b8cee) * $signed(16'h1);
  assign T10392 = T10390[6'h2d:6'h2d];
  assign T10393 = T2943[1'h0:1'h0];
  assign T10394 = T10407 ? twiddle4_3_467_real : twiddle4_3_466_real;
  assign twiddle4_3_466_real = T10397 + T10395;
  assign T10395 = $signed(T10396) / $signed(22'h100000);
  assign T10396 = $signed(31'h45a69bbf) * $signed(16'h0);
  assign T10397 = {T10400, T10398};
  assign T10398 = $signed(T10399) / $signed(22'h100000);
  assign T10399 = $signed(30'h25b4bed9) * $signed(16'h1);
  assign T10400 = T10398[6'h2d:6'h2d];
  assign twiddle4_3_467_real = T10403 + T10401;
  assign T10401 = $signed(T10402) / $signed(22'h100000);
  assign T10402 = $signed(31'h456949ca) * $signed(16'h0);
  assign T10403 = {T10406, T10404};
  assign T10404 = $signed(T10405) / $signed(22'h100000);
  assign T10405 = $signed(30'h263e82bc) * $signed(16'h1);
  assign T10406 = T10404[6'h2d:6'h2d];
  assign T10407 = T2943[1'h0:1'h0];
  assign T10408 = T2943[1'h1:1'h1];
  assign T10409 = T10438 ? T10424 : T10410;
  assign T10410 = T10423 ? twiddle4_3_469_real : twiddle4_3_468_real;
  assign twiddle4_3_468_real = T10413 + T10411;
  assign T10411 = $signed(T10412) / $signed(22'h100000);
  assign T10412 = $signed(31'h452d3d19) * $signed(16'h0);
  assign T10413 = {T10416, T10414};
  assign T10414 = $signed(T10415) / $signed(22'h100000);
  assign T10415 = $signed(30'h26c8d59d) * $signed(16'h1);
  assign T10416 = T10414[6'h2d:6'h2d];
  assign twiddle4_3_469_real = T10419 + T10417;
  assign T10417 = $signed(T10418) / $signed(22'h100000);
  assign T10418 = $signed(31'h44f276f8) * $signed(16'h0);
  assign T10419 = {T10422, T10420};
  assign T10420 = $signed(T10421) / $signed(22'h100000);
  assign T10421 = $signed(30'h2753b47a) * $signed(16'h1);
  assign T10422 = T10420[6'h2d:6'h2d];
  assign T10423 = T2943[1'h0:1'h0];
  assign T10424 = T10437 ? twiddle4_3_471_real : twiddle4_3_470_real;
  assign twiddle4_3_470_real = T10427 + T10425;
  assign T10425 = $signed(T10426) / $signed(22'h100000);
  assign T10426 = $signed(31'h44b8f8ae) * $signed(16'h0);
  assign T10427 = {T10430, T10428};
  assign T10428 = $signed(T10429) / $signed(22'h100000);
  assign T10429 = $signed(30'h27df1c50) * $signed(16'h1);
  assign T10430 = T10428[6'h2d:6'h2d];
  assign twiddle4_3_471_real = T10433 + T10431;
  assign T10431 = $signed(T10432) / $signed(22'h100000);
  assign T10432 = $signed(31'h4480c379) * $signed(16'h0);
  assign T10433 = {T10436, T10434};
  assign T10434 = $signed(T10435) / $signed(22'h100000);
  assign T10435 = $signed(30'h286b0a1a) * $signed(16'h1);
  assign T10436 = T10434[6'h2d:6'h2d];
  assign T10437 = T2943[1'h0:1'h0];
  assign T10438 = T2943[1'h1:1'h1];
  assign T10439 = T2943[2'h2:2'h2];
  assign T10440 = T10501 ? T10471 : T10441;
  assign T10441 = T10470 ? T10456 : T10442;
  assign T10442 = T10455 ? twiddle4_3_473_real : twiddle4_3_472_real;
  assign twiddle4_3_472_real = T10445 + T10443;
  assign T10443 = $signed(T10444) / $signed(22'h100000);
  assign T10444 = $signed(31'h4449d893) * $signed(16'h0);
  assign T10445 = {T10448, T10446};
  assign T10446 = $signed(T10447) / $signed(22'h100000);
  assign T10447 = $signed(30'h28f77ad0) * $signed(16'h1);
  assign T10448 = T10446[6'h2d:6'h2d];
  assign twiddle4_3_473_real = T10451 + T10449;
  assign T10449 = $signed(T10450) / $signed(22'h100000);
  assign T10450 = $signed(31'h4414392b) * $signed(16'h0);
  assign T10451 = {T10454, T10452};
  assign T10452 = $signed(T10453) / $signed(22'h100000);
  assign T10453 = $signed(30'h29846b64) * $signed(16'h1);
  assign T10454 = T10452[6'h2d:6'h2d];
  assign T10455 = T2943[1'h0:1'h0];
  assign T10456 = T10469 ? twiddle4_3_475_real : twiddle4_3_474_real;
  assign twiddle4_3_474_real = T10459 + T10457;
  assign T10457 = $signed(T10458) / $signed(22'h100000);
  assign T10458 = $signed(31'h43dfe66c) * $signed(16'h0);
  assign T10459 = {T10462, T10460};
  assign T10460 = $signed(T10461) / $signed(22'h100000);
  assign T10461 = $signed(30'h2a11d8c9) * $signed(16'h1);
  assign T10462 = T10460[6'h2d:6'h2d];
  assign twiddle4_3_475_real = T10465 + T10463;
  assign T10463 = $signed(T10464) / $signed(22'h100000);
  assign T10464 = $signed(31'h43ace178) * $signed(16'h0);
  assign T10465 = {T10468, T10466};
  assign T10466 = $signed(T10467) / $signed(22'h100000);
  assign T10467 = $signed(30'h2a9fbfee) * $signed(16'h1);
  assign T10468 = T10466[6'h2d:6'h2d];
  assign T10469 = T2943[1'h0:1'h0];
  assign T10470 = T2943[1'h1:1'h1];
  assign T10471 = T10500 ? T10486 : T10472;
  assign T10472 = T10485 ? twiddle4_3_477_real : twiddle4_3_476_real;
  assign twiddle4_3_476_real = T10475 + T10473;
  assign T10473 = $signed(T10474) / $signed(22'h100000);
  assign T10474 = $signed(31'h437b2b6a) * $signed(16'h0);
  assign T10475 = {T10478, T10476};
  assign T10476 = $signed(T10477) / $signed(22'h100000);
  assign T10477 = $signed(30'h2b2e1dbe) * $signed(16'h1);
  assign T10478 = T10476[6'h2d:6'h2d];
  assign twiddle4_3_477_real = T10481 + T10479;
  assign T10479 = $signed(T10480) / $signed(22'h100000);
  assign T10480 = $signed(31'h434ac556) * $signed(16'h0);
  assign T10481 = {T10484, T10482};
  assign T10482 = $signed(T10483) / $signed(22'h100000);
  assign T10483 = $signed(30'h2bbcef24) * $signed(16'h1);
  assign T10484 = T10482[6'h2d:6'h2d];
  assign T10485 = T2943[1'h0:1'h0];
  assign T10486 = T10499 ? twiddle4_3_479_real : twiddle4_3_478_real;
  assign twiddle4_3_478_real = T10489 + T10487;
  assign T10487 = $signed(T10488) / $signed(22'h100000);
  assign T10488 = $signed(31'h431bb04a) * $signed(16'h0);
  assign T10489 = {T10492, T10490};
  assign T10490 = $signed(T10491) / $signed(22'h100000);
  assign T10491 = $signed(30'h2c4c3106) * $signed(16'h1);
  assign T10492 = T10490[6'h2d:6'h2d];
  assign twiddle4_3_479_real = T10495 + T10493;
  assign T10493 = $signed(T10494) / $signed(22'h100000);
  assign T10494 = $signed(31'h42eded49) * $signed(16'h0);
  assign T10495 = {T10498, T10496};
  assign T10496 = $signed(T10497) / $signed(22'h100000);
  assign T10497 = $signed(30'h2cdbe04a) * $signed(16'h1);
  assign T10498 = T10496[6'h2d:6'h2d];
  assign T10499 = T2943[1'h0:1'h0];
  assign T10500 = T2943[1'h1:1'h1];
  assign T10501 = T2943[2'h2:2'h2];
  assign T10502 = T2943[2'h3:2'h3];
  assign T10503 = T2943[3'h4:3'h4];
  assign T10504 = T10784 ? T10642 : T10505;
  assign T10505 = T10641 ? T10571 : T10506;
  assign T10506 = T10570 ? T10537 : T10507;
  assign T10507 = T10536 ? T10522 : T10508;
  assign T10508 = T10521 ? twiddle4_3_481_real : twiddle4_3_480_real;
  assign twiddle4_3_480_real = T10511 + T10509;
  assign T10509 = $signed(T10510) / $signed(22'h100000);
  assign T10510 = $signed(31'h42c17d53) * $signed(16'h0);
  assign T10511 = {T10514, T10512};
  assign T10512 = $signed(T10513) / $signed(22'h100000);
  assign T10513 = $signed(30'h2d6bf9d2) * $signed(16'h1);
  assign T10514 = T10512[6'h2d:6'h2d];
  assign twiddle4_3_481_real = T10517 + T10515;
  assign T10515 = $signed(T10516) / $signed(22'h100000);
  assign T10516 = $signed(31'h4296615e) * $signed(16'h0);
  assign T10517 = {T10520, T10518};
  assign T10518 = $signed(T10519) / $signed(22'h100000);
  assign T10519 = $signed(30'h2dfc7a7d) * $signed(16'h1);
  assign T10520 = T10518[6'h2d:6'h2d];
  assign T10521 = T2943[1'h0:1'h0];
  assign T10522 = T10535 ? twiddle4_3_483_real : twiddle4_3_482_real;
  assign twiddle4_3_482_real = T10525 + T10523;
  assign T10523 = $signed(T10524) / $signed(22'h100000);
  assign T10524 = $signed(31'h426c9a59) * $signed(16'h0);
  assign T10525 = {T10528, T10526};
  assign T10526 = $signed(T10527) / $signed(22'h100000);
  assign T10527 = $signed(30'h2e8d5f29) * $signed(16'h1);
  assign T10528 = T10526[6'h2d:6'h2d];
  assign twiddle4_3_483_real = T10531 + T10529;
  assign T10529 = $signed(T10530) / $signed(22'h100000);
  assign T10530 = $signed(31'h4244292c) * $signed(16'h0);
  assign T10531 = {T10534, T10532};
  assign T10532 = $signed(T10533) / $signed(22'h100000);
  assign T10533 = $signed(30'h2f1ea4b2) * $signed(16'h1);
  assign T10534 = T10532[6'h2d:6'h2d];
  assign T10535 = T2943[1'h0:1'h0];
  assign T10536 = T2943[1'h1:1'h1];
  assign T10537 = T10569 ? T10553 : T10538;
  assign T10538 = T10552 ? twiddle4_3_485_real : twiddle4_3_484_real;
  assign twiddle4_3_484_real = T10541 + T10539;
  assign T10539 = $signed(T10540) / $signed(22'h100000);
  assign T10540 = $signed(31'h421d0eb9) * $signed(16'h0);
  assign T10541 = {T10544, T10542};
  assign T10542 = $signed(T10543) / $signed(22'h100000);
  assign T10543 = $signed(30'h2fb047f2) * $signed(16'h1);
  assign T10544 = T10542[6'h2d:6'h2d];
  assign twiddle4_3_485_real = T10547 + T10545;
  assign T10545 = $signed(T10546) / $signed(22'h100000);
  assign T10546 = $signed(31'h41f74bd7) * $signed(16'h0);
  assign T10547 = {T10550, T10548};
  assign T10548 = $signed(T10549) / $signed(22'h100000);
  assign T10549 = $signed(29'h104245c0) * $signed(16'h1);
  assign T10550 = T10551 ? 2'h3 : 2'h0;
  assign T10551 = T10548[6'h2c:6'h2c];
  assign T10552 = T2943[1'h0:1'h0];
  assign T10553 = T10568 ? twiddle4_3_487_real : twiddle4_3_486_real;
  assign twiddle4_3_486_real = T10556 + T10554;
  assign T10554 = $signed(T10555) / $signed(22'h100000);
  assign T10555 = $signed(31'h41d2e159) * $signed(16'h0);
  assign T10556 = {T10559, T10557};
  assign T10557 = $signed(T10558) / $signed(22'h100000);
  assign T10558 = $signed(29'h10d49af1) * $signed(16'h1);
  assign T10559 = T10560 ? 2'h3 : 2'h0;
  assign T10560 = T10557[6'h2c:6'h2c];
  assign twiddle4_3_487_real = T10563 + T10561;
  assign T10561 = $signed(T10562) / $signed(22'h100000);
  assign T10562 = $signed(31'h41afd008) * $signed(16'h0);
  assign T10563 = {T10566, T10564};
  assign T10564 = $signed(T10565) / $signed(22'h100000);
  assign T10565 = $signed(29'h1167445a) * $signed(16'h1);
  assign T10566 = T10567 ? 2'h3 : 2'h0;
  assign T10567 = T10564[6'h2c:6'h2c];
  assign T10568 = T2943[1'h0:1'h0];
  assign T10569 = T2943[1'h1:1'h1];
  assign T10570 = T2943[2'h2:2'h2];
  assign T10571 = T10640 ? T10606 : T10572;
  assign T10572 = T10605 ? T10589 : T10573;
  assign T10573 = T10588 ? twiddle4_3_489_real : twiddle4_3_488_real;
  assign twiddle4_3_488_real = T10576 + T10574;
  assign T10574 = $signed(T10575) / $signed(22'h100000);
  assign T10575 = $signed(31'h418e18a8) * $signed(16'h0);
  assign T10576 = {T10579, T10577};
  assign T10577 = $signed(T10578) / $signed(22'h100000);
  assign T10578 = $signed(29'h11fa3ecb) * $signed(16'h1);
  assign T10579 = T10580 ? 2'h3 : 2'h0;
  assign T10580 = T10577[6'h2c:6'h2c];
  assign twiddle4_3_489_real = T10583 + T10581;
  assign T10581 = $signed(T10582) / $signed(22'h100000);
  assign T10582 = $signed(31'h416dbbf3) * $signed(16'h0);
  assign T10583 = {T10586, T10584};
  assign T10584 = $signed(T10585) / $signed(22'h100000);
  assign T10585 = $signed(29'h128d8716) * $signed(16'h1);
  assign T10586 = T10587 ? 2'h3 : 2'h0;
  assign T10587 = T10584[6'h2c:6'h2c];
  assign T10588 = T2943[1'h0:1'h0];
  assign T10589 = T10604 ? twiddle4_3_491_real : twiddle4_3_490_real;
  assign twiddle4_3_490_real = T10592 + T10590;
  assign T10590 = $signed(T10591) / $signed(22'h100000);
  assign T10591 = $signed(31'h414eba9e) * $signed(16'h0);
  assign T10592 = {T10595, T10593};
  assign T10593 = $signed(T10594) / $signed(22'h100000);
  assign T10594 = $signed(29'h13211a07) * $signed(16'h1);
  assign T10595 = T10596 ? 2'h3 : 2'h0;
  assign T10596 = T10593[6'h2c:6'h2c];
  assign twiddle4_3_491_real = T10599 + T10597;
  assign T10597 = $signed(T10598) / $signed(22'h100000);
  assign T10598 = $signed(31'h41311553) * $signed(16'h0);
  assign T10599 = {T10602, T10600};
  assign T10600 = $signed(T10601) / $signed(22'h100000);
  assign T10601 = $signed(29'h13b4f46d) * $signed(16'h1);
  assign T10602 = T10603 ? 2'h3 : 2'h0;
  assign T10603 = T10600[6'h2c:6'h2c];
  assign T10604 = T2943[1'h0:1'h0];
  assign T10605 = T2943[1'h1:1'h1];
  assign T10606 = T10639 ? T10623 : T10607;
  assign T10607 = T10622 ? twiddle4_3_493_real : twiddle4_3_492_real;
  assign twiddle4_3_492_real = T10610 + T10608;
  assign T10608 = $signed(T10609) / $signed(22'h100000);
  assign T10609 = $signed(31'h4114ccb9) * $signed(16'h0);
  assign T10610 = {T10613, T10611};
  assign T10611 = $signed(T10612) / $signed(22'h100000);
  assign T10612 = $signed(29'h14491311) * $signed(16'h1);
  assign T10613 = T10614 ? 2'h3 : 2'h0;
  assign T10614 = T10611[6'h2c:6'h2c];
  assign twiddle4_3_493_real = T10617 + T10615;
  assign T10615 = $signed(T10616) / $signed(22'h100000);
  assign T10616 = $signed(31'h40f9e16c) * $signed(16'h0);
  assign T10617 = {T10620, T10618};
  assign T10618 = $signed(T10619) / $signed(22'h100000);
  assign T10619 = $signed(29'h14dd72bf) * $signed(16'h1);
  assign T10620 = T10621 ? 2'h3 : 2'h0;
  assign T10621 = T10618[6'h2c:6'h2c];
  assign T10622 = T2943[1'h0:1'h0];
  assign T10623 = T10638 ? twiddle4_3_495_real : twiddle4_3_494_real;
  assign twiddle4_3_494_real = T10626 + T10624;
  assign T10624 = $signed(T10625) / $signed(22'h100000);
  assign T10625 = $signed(31'h40e05401) * $signed(16'h0);
  assign T10626 = {T10629, T10627};
  assign T10627 = $signed(T10628) / $signed(22'h100000);
  assign T10628 = $signed(29'h1572103e) * $signed(16'h1);
  assign T10629 = T10630 ? 2'h3 : 2'h0;
  assign T10630 = T10627[6'h2c:6'h2c];
  assign twiddle4_3_495_real = T10633 + T10631;
  assign T10631 = $signed(T10632) / $signed(22'h100000);
  assign T10632 = $signed(31'h40c82507) * $signed(16'h0);
  assign T10633 = {T10636, T10634};
  assign T10634 = $signed(T10635) / $signed(22'h100000);
  assign T10635 = $signed(29'h1606e855) * $signed(16'h1);
  assign T10636 = T10637 ? 2'h3 : 2'h0;
  assign T10637 = T10634[6'h2c:6'h2c];
  assign T10638 = T2943[1'h0:1'h0];
  assign T10639 = T2943[1'h1:1'h1];
  assign T10640 = T2943[2'h2:2'h2];
  assign T10641 = T2943[2'h3:2'h3];
  assign T10642 = T10783 ? T10713 : T10643;
  assign T10643 = T10712 ? T10678 : T10644;
  assign T10644 = T10677 ? T10661 : T10645;
  assign T10645 = T10660 ? twiddle4_3_497_real : twiddle4_3_496_real;
  assign twiddle4_3_496_real = T10648 + T10646;
  assign T10646 = $signed(T10647) / $signed(22'h100000);
  assign T10647 = $signed(31'h40b15502) * $signed(16'h0);
  assign T10648 = {T10651, T10649};
  assign T10649 = $signed(T10650) / $signed(22'h100000);
  assign T10650 = $signed(29'h169bf7c9) * $signed(16'h1);
  assign T10651 = T10652 ? 2'h3 : 2'h0;
  assign T10652 = T10649[6'h2c:6'h2c];
  assign twiddle4_3_497_real = T10655 + T10653;
  assign T10653 = $signed(T10654) / $signed(22'h100000);
  assign T10654 = $signed(31'h409be473) * $signed(16'h0);
  assign T10655 = {T10658, T10656};
  assign T10656 = $signed(T10657) / $signed(22'h100000);
  assign T10657 = $signed(29'h17313b60) * $signed(16'h1);
  assign T10658 = T10659 ? 2'h3 : 2'h0;
  assign T10659 = T10656[6'h2c:6'h2c];
  assign T10660 = T2943[1'h0:1'h0];
  assign T10661 = T10676 ? twiddle4_3_499_real : twiddle4_3_498_real;
  assign twiddle4_3_498_real = T10664 + T10662;
  assign T10662 = $signed(T10663) / $signed(22'h100000);
  assign T10663 = $signed(31'h4087d3d1) * $signed(16'h0);
  assign T10664 = {T10667, T10665};
  assign T10665 = $signed(T10666) / $signed(22'h100000);
  assign T10666 = $signed(29'h17c6afdd) * $signed(16'h1);
  assign T10667 = T10668 ? 2'h3 : 2'h0;
  assign T10668 = T10665[6'h2c:6'h2c];
  assign twiddle4_3_499_real = T10671 + T10669;
  assign T10669 = $signed(T10670) / $signed(22'h100000);
  assign T10670 = $signed(31'h4075238a) * $signed(16'h0);
  assign T10671 = {T10674, T10672};
  assign T10672 = $signed(T10673) / $signed(22'h100000);
  assign T10673 = $signed(28'h85c5201) * $signed(16'h1);
  assign T10674 = T10675 ? 3'h7 : 3'h0;
  assign T10675 = T10672[6'h2b:6'h2b];
  assign T10676 = T2943[1'h0:1'h0];
  assign T10677 = T2943[1'h1:1'h1];
  assign T10678 = T10711 ? T10695 : T10679;
  assign T10679 = T10694 ? twiddle4_3_501_real : twiddle4_3_500_real;
  assign twiddle4_3_500_real = T10682 + T10680;
  assign T10680 = $signed(T10681) / $signed(22'h100000);
  assign T10681 = $signed(31'h4063d406) * $signed(16'h0);
  assign T10682 = {T10685, T10683};
  assign T10683 = $signed(T10684) / $signed(22'h100000);
  assign T10684 = $signed(28'h8f21e8f) * $signed(16'h1);
  assign T10685 = T10686 ? 3'h7 : 3'h0;
  assign T10686 = T10683[6'h2b:6'h2b];
  assign twiddle4_3_501_real = T10689 + T10687;
  assign T10687 = $signed(T10688) / $signed(22'h100000);
  assign T10688 = $signed(31'h4053e5a5) * $signed(16'h0);
  assign T10689 = {T10692, T10690};
  assign T10690 = $signed(T10691) / $signed(22'h100000);
  assign T10691 = $signed(28'h9881246) * $signed(16'h1);
  assign T10692 = T10693 ? 3'h7 : 3'h0;
  assign T10693 = T10690[6'h2b:6'h2b];
  assign T10694 = T2943[1'h0:1'h0];
  assign T10695 = T10710 ? twiddle4_3_503_real : twiddle4_3_502_real;
  assign twiddle4_3_502_real = T10698 + T10696;
  assign T10696 = $signed(T10697) / $signed(22'h100000);
  assign T10697 = $signed(31'h404558c1) * $signed(16'h0);
  assign T10698 = {T10701, T10699};
  assign T10699 = $signed(T10700) / $signed(22'h100000);
  assign T10700 = $signed(28'ha1e29e6) * $signed(16'h1);
  assign T10701 = T10702 ? 3'h7 : 3'h0;
  assign T10702 = T10699[6'h2b:6'h2b];
  assign twiddle4_3_503_real = T10705 + T10703;
  assign T10703 = $signed(T10704) / $signed(22'h100000);
  assign T10704 = $signed(31'h40382da9) * $signed(16'h0);
  assign T10705 = {T10708, T10706};
  assign T10706 = $signed(T10707) / $signed(22'h100000);
  assign T10707 = $signed(28'hab4622e) * $signed(16'h1);
  assign T10708 = T10709 ? 3'h7 : 3'h0;
  assign T10709 = T10706[6'h2b:6'h2b];
  assign T10710 = T2943[1'h0:1'h0];
  assign T10711 = T2943[1'h1:1'h1];
  assign T10712 = T2943[2'h2:2'h2];
  assign T10713 = T10782 ? T10748 : T10714;
  assign T10714 = T10747 ? T10731 : T10715;
  assign T10715 = T10730 ? twiddle4_3_505_real : twiddle4_3_504_real;
  assign twiddle4_3_504_real = T10718 + T10716;
  assign T10716 = $signed(T10717) / $signed(22'h100000);
  assign T10717 = $signed(31'h402c64a6) * $signed(16'h0);
  assign T10718 = {T10721, T10719};
  assign T10719 = $signed(T10720) / $signed(22'h100000);
  assign T10720 = $signed(28'hb4ab7dc) * $signed(16'h1);
  assign T10721 = T10722 ? 3'h7 : 3'h0;
  assign T10722 = T10719[6'h2b:6'h2b];
  assign twiddle4_3_505_real = T10725 + T10723;
  assign T10723 = $signed(T10724) / $signed(22'h100000);
  assign T10724 = $signed(31'h4021fdfb) * $signed(16'h0);
  assign T10725 = {T10728, T10726};
  assign T10726 = $signed(T10727) / $signed(22'h100000);
  assign T10727 = $signed(28'hbe127ad) * $signed(16'h1);
  assign T10728 = T10729 ? 3'h7 : 3'h0;
  assign T10729 = T10726[6'h2b:6'h2b];
  assign T10730 = T2943[1'h0:1'h0];
  assign T10731 = T10746 ? twiddle4_3_507_real : twiddle4_3_506_real;
  assign twiddle4_3_506_real = T10734 + T10732;
  assign T10732 = $signed(T10733) / $signed(22'h100000);
  assign T10733 = $signed(31'h4018f9e1) * $signed(16'h0);
  assign T10734 = {T10737, T10735};
  assign T10735 = $signed(T10736) / $signed(22'h100000);
  assign T10736 = $signed(27'h477ae5e) * $signed(16'h1);
  assign T10737 = T10738 ? 4'hf : 4'h0;
  assign T10738 = T10735[6'h2a:6'h2a];
  assign twiddle4_3_507_real = T10741 + T10739;
  assign T10739 = $signed(T10740) / $signed(22'h100000);
  assign T10740 = $signed(31'h4011588a) * $signed(16'h0);
  assign T10741 = {T10744, T10742};
  assign T10742 = $signed(T10743) / $signed(22'h100000);
  assign T10743 = $signed(27'h50e48ac) * $signed(16'h1);
  assign T10744 = T10745 ? 4'hf : 4'h0;
  assign T10745 = T10742[6'h2a:6'h2a];
  assign T10746 = T2943[1'h0:1'h0];
  assign T10747 = T2943[1'h1:1'h1];
  assign T10748 = T10781 ? T10765 : T10749;
  assign T10749 = T10764 ? twiddle4_3_509_real : twiddle4_3_508_real;
  assign twiddle4_3_508_real = T10752 + T10750;
  assign T10750 = $signed(T10751) / $signed(22'h100000);
  assign T10751 = $signed(31'h400b1a21) * $signed(16'h0);
  assign T10752 = {T10755, T10753};
  assign T10753 = $signed(T10754) / $signed(22'h100000);
  assign T10754 = $signed(27'h5a4f352) * $signed(16'h1);
  assign T10755 = T10756 ? 4'hf : 4'h0;
  assign T10756 = T10753[6'h2a:6'h2a];
  assign twiddle4_3_509_real = T10759 + T10757;
  assign T10757 = $signed(T10758) / $signed(22'h100000);
  assign T10758 = $signed(31'h40063ec7) * $signed(16'h0);
  assign T10759 = {T10762, T10760};
  assign T10760 = $signed(T10761) / $signed(22'h100000);
  assign T10761 = $signed(26'h23bab0c) * $signed(16'h1);
  assign T10762 = T10763 ? 5'h1f : 5'h0;
  assign T10763 = T10760[6'h29:6'h29];
  assign T10764 = T2943[1'h0:1'h0];
  assign T10765 = T10780 ? twiddle4_3_511_real : twiddle4_3_510_real;
  assign twiddle4_3_510_real = T10768 + T10766;
  assign T10766 = $signed(T10767) / $signed(22'h100000);
  assign T10767 = $signed(31'h4002c698) * $signed(16'h0);
  assign T10768 = {T10771, T10769};
  assign T10769 = $signed(T10770) / $signed(22'h100000);
  assign T10770 = $signed(26'h2d26c95) * $signed(16'h1);
  assign T10771 = T10772 ? 5'h1f : 5'h0;
  assign T10772 = T10769[6'h29:6'h29];
  assign twiddle4_3_511_real = T10775 + T10773;
  assign T10773 = $signed(T10774) / $signed(22'h100000);
  assign T10774 = $signed(31'h4000b1a7) * $signed(16'h0);
  assign T10775 = {T10778, T10776};
  assign T10776 = $signed(T10777) / $signed(22'h100000);
  assign T10777 = $signed(25'h16934a8) * $signed(16'h1);
  assign T10778 = T10779 ? 6'h3f : 6'h0;
  assign T10779 = T10776[6'h28:6'h28];
  assign T10780 = T2943[1'h0:1'h0];
  assign T10781 = T2943[1'h1:1'h1];
  assign T10782 = T2943[2'h2:2'h2];
  assign T10783 = T2943[2'h3:2'h3];
  assign T10784 = T2943[3'h4:3'h4];
  assign T10785 = T2943[3'h5:3'h5];
  assign T10786 = T2943[3'h6:3'h6];
  assign T10787 = T2943[3'h7:3'h7];
  assign T10788 = T8832[6'h2e:6'h2e];
  assign T10789 = T2943[4'h8:4'h8];
  assign io_t4_2out_imag = T10790;
  assign T10790 = T10791[4'hf:1'h0];
  assign T10791 = T14744 ? T12769 : T10792;
  assign T10792 = T12768 ? T11789 : T10793;
  assign T10793 = T11788 ? T11360 : T10794;
  assign T10794 = T11359 ? T11093 : T10795;
  assign T10795 = T11092 ? T10948 : T10796;
  assign T10796 = T10947 ? T10875 : T10797;
  assign T10797 = T10874 ? T10838 : T10798;
  assign T10798 = T10837 ? T10819 : T10799;
  assign T10799 = T10816 ? T10807 : twiddle4_2_0_imag;
  assign twiddle4_2_0_imag = T10805 + T10800;
  assign T10800 = {T10803, T10801};
  assign T10801 = $signed(T10802) / $signed(22'h100000);
  assign T10802 = $signed(1'h0) * $signed(16'hffff);
  assign T10803 = T10804 ? 31'h7fffffff : 31'h0;
  assign T10804 = T10801[5'h10:5'h10];
  assign T10805 = $signed(T10806) / $signed(22'h100000);
  assign T10806 = $signed(32'h40000000) * $signed(16'h0);
  assign T10807 = {T10815, twiddle4_2_1_imag};
  assign twiddle4_2_1_imag = T10813 + T10808;
  assign T10808 = {T10811, T10809};
  assign T10809 = $signed(T10810) / $signed(22'h100000);
  assign T10810 = $signed(24'h6487c3) * $signed(16'hffff);
  assign T10811 = T10812 ? 7'h7f : 7'h0;
  assign T10812 = T10809[6'h27:6'h27];
  assign T10813 = $signed(T10814) / $signed(22'h100000);
  assign T10814 = $signed(31'h3fffb10b) * $signed(16'h0);
  assign T10815 = twiddle4_2_1_imag[6'h2e:6'h2e];
  assign T10816 = T10817[1'h0:1'h0];
  assign T10817 = T10818;
  assign T10818 = io_in4[4'h8:1'h0];
  assign T10819 = {T10836, T10820};
  assign T10820 = T10835 ? twiddle4_2_3_imag : twiddle4_2_2_imag;
  assign twiddle4_2_2_imag = T10826 + T10821;
  assign T10821 = {T10824, T10822};
  assign T10822 = $signed(T10823) / $signed(22'h100000);
  assign T10823 = $signed(25'hc90e8f) * $signed(16'hffff);
  assign T10824 = T10825 ? 6'h3f : 6'h0;
  assign T10825 = T10822[6'h28:6'h28];
  assign T10826 = $signed(T10827) / $signed(22'h100000);
  assign T10827 = $signed(31'h3ffec42d) * $signed(16'h0);
  assign twiddle4_2_3_imag = T10833 + T10828;
  assign T10828 = {T10831, T10829};
  assign T10829 = $signed(T10830) / $signed(22'h100000);
  assign T10830 = $signed(26'h12d936b) * $signed(16'hffff);
  assign T10831 = T10832 ? 5'h1f : 5'h0;
  assign T10832 = T10829[6'h29:6'h29];
  assign T10833 = $signed(T10834) / $signed(22'h100000);
  assign T10834 = $signed(31'h3ffd3968) * $signed(16'h0);
  assign T10835 = T10817[1'h0:1'h0];
  assign T10836 = T10820[6'h2e:6'h2e];
  assign T10837 = T10817[1'h1:1'h1];
  assign T10838 = {T10873, T10839};
  assign T10839 = T10872 ? T10856 : T10840;
  assign T10840 = T10855 ? twiddle4_2_5_imag : twiddle4_2_4_imag;
  assign twiddle4_2_4_imag = T10846 + T10841;
  assign T10841 = {T10844, T10842};
  assign T10842 = $signed(T10843) / $signed(22'h100000);
  assign T10843 = $signed(26'h192155f) * $signed(16'hffff);
  assign T10844 = T10845 ? 5'h1f : 5'h0;
  assign T10845 = T10842[6'h29:6'h29];
  assign T10846 = $signed(T10847) / $signed(22'h100000);
  assign T10847 = $signed(31'h3ffb10c1) * $signed(16'h0);
  assign twiddle4_2_5_imag = T10853 + T10848;
  assign T10848 = {T10851, T10849};
  assign T10849 = $signed(T10850) / $signed(22'h100000);
  assign T10850 = $signed(26'h1f69373) * $signed(16'hffff);
  assign T10851 = T10852 ? 5'h1f : 5'h0;
  assign T10852 = T10849[6'h29:6'h29];
  assign T10853 = $signed(T10854) / $signed(22'h100000);
  assign T10854 = $signed(31'h3ff84a3b) * $signed(16'h0);
  assign T10855 = T10817[1'h0:1'h0];
  assign T10856 = T10871 ? twiddle4_2_7_imag : twiddle4_2_6_imag;
  assign twiddle4_2_6_imag = T10862 + T10857;
  assign T10857 = {T10860, T10858};
  assign T10858 = $signed(T10859) / $signed(22'h100000);
  assign T10859 = $signed(27'h25b0cae) * $signed(16'hffff);
  assign T10860 = T10861 ? 4'hf : 4'h0;
  assign T10861 = T10858[6'h2a:6'h2a];
  assign T10862 = $signed(T10863) / $signed(22'h100000);
  assign T10863 = $signed(31'h3ff4e5df) * $signed(16'h0);
  assign twiddle4_2_7_imag = T10869 + T10864;
  assign T10864 = {T10867, T10865};
  assign T10865 = $signed(T10866) / $signed(22'h100000);
  assign T10866 = $signed(27'h2bf801a) * $signed(16'hffff);
  assign T10867 = T10868 ? 4'hf : 4'h0;
  assign T10868 = T10865[6'h2a:6'h2a];
  assign T10869 = $signed(T10870) / $signed(22'h100000);
  assign T10870 = $signed(31'h3ff0e3b5) * $signed(16'h0);
  assign T10871 = T10817[1'h0:1'h0];
  assign T10872 = T10817[1'h1:1'h1];
  assign T10873 = T10839[6'h2e:6'h2e];
  assign T10874 = T10817[2'h2:2'h2];
  assign T10875 = {T10946, T10876};
  assign T10876 = T10945 ? T10911 : T10877;
  assign T10877 = T10910 ? T10894 : T10878;
  assign T10878 = T10893 ? twiddle4_2_9_imag : twiddle4_2_8_imag;
  assign twiddle4_2_8_imag = T10884 + T10879;
  assign T10879 = {T10882, T10880};
  assign T10880 = $signed(T10881) / $signed(22'h100000);
  assign T10881 = $signed(27'h323ecbe) * $signed(16'hffff);
  assign T10882 = T10883 ? 4'hf : 4'h0;
  assign T10883 = T10880[6'h2a:6'h2a];
  assign T10884 = $signed(T10885) / $signed(22'h100000);
  assign T10885 = $signed(31'h3fec43c6) * $signed(16'h0);
  assign twiddle4_2_9_imag = T10891 + T10886;
  assign T10886 = {T10889, T10887};
  assign T10887 = $signed(T10888) / $signed(22'h100000);
  assign T10888 = $signed(27'h38851a2) * $signed(16'hffff);
  assign T10889 = T10890 ? 4'hf : 4'h0;
  assign T10890 = T10887[6'h2a:6'h2a];
  assign T10891 = $signed(T10892) / $signed(22'h100000);
  assign T10892 = $signed(31'h3fe7061f) * $signed(16'h0);
  assign T10893 = T10817[1'h0:1'h0];
  assign T10894 = T10909 ? twiddle4_2_11_imag : twiddle4_2_10_imag;
  assign twiddle4_2_10_imag = T10900 + T10895;
  assign T10895 = {T10898, T10896};
  assign T10896 = $signed(T10897) / $signed(22'h100000);
  assign T10897 = $signed(27'h3ecadcf) * $signed(16'hffff);
  assign T10898 = T10899 ? 4'hf : 4'h0;
  assign T10899 = T10896[6'h2a:6'h2a];
  assign T10900 = $signed(T10901) / $signed(22'h100000);
  assign T10901 = $signed(31'h3fe12acb) * $signed(16'h0);
  assign twiddle4_2_11_imag = T10907 + T10902;
  assign T10902 = {T10905, T10903};
  assign T10903 = $signed(T10904) / $signed(22'h100000);
  assign T10904 = $signed(28'h451004d) * $signed(16'hffff);
  assign T10905 = T10906 ? 3'h7 : 3'h0;
  assign T10906 = T10903[6'h2b:6'h2b];
  assign T10907 = $signed(T10908) / $signed(22'h100000);
  assign T10908 = $signed(31'h3fdab1d9) * $signed(16'h0);
  assign T10909 = T10817[1'h0:1'h0];
  assign T10910 = T10817[1'h1:1'h1];
  assign T10911 = T10944 ? T10928 : T10912;
  assign T10912 = T10927 ? twiddle4_2_13_imag : twiddle4_2_12_imag;
  assign twiddle4_2_12_imag = T10918 + T10913;
  assign T10913 = {T10916, T10914};
  assign T10914 = $signed(T10915) / $signed(22'h100000);
  assign T10915 = $signed(28'h4b54824) * $signed(16'hffff);
  assign T10916 = T10917 ? 3'h7 : 3'h0;
  assign T10917 = T10914[6'h2b:6'h2b];
  assign T10918 = $signed(T10919) / $signed(22'h100000);
  assign T10919 = $signed(31'h3fd39b5a) * $signed(16'h0);
  assign twiddle4_2_13_imag = T10925 + T10920;
  assign T10920 = {T10923, T10921};
  assign T10921 = $signed(T10922) / $signed(22'h100000);
  assign T10922 = $signed(28'h519845e) * $signed(16'hffff);
  assign T10923 = T10924 ? 3'h7 : 3'h0;
  assign T10924 = T10921[6'h2b:6'h2b];
  assign T10925 = $signed(T10926) / $signed(22'h100000);
  assign T10926 = $signed(31'h3fcbe75e) * $signed(16'h0);
  assign T10927 = T10817[1'h0:1'h0];
  assign T10928 = T10943 ? twiddle4_2_15_imag : twiddle4_2_14_imag;
  assign twiddle4_2_14_imag = T10934 + T10929;
  assign T10929 = {T10932, T10930};
  assign T10930 = $signed(T10931) / $signed(22'h100000);
  assign T10931 = $signed(28'h57db402) * $signed(16'hffff);
  assign T10932 = T10933 ? 3'h7 : 3'h0;
  assign T10933 = T10930[6'h2b:6'h2b];
  assign T10934 = $signed(T10935) / $signed(22'h100000);
  assign T10935 = $signed(31'h3fc395f9) * $signed(16'h0);
  assign twiddle4_2_15_imag = T10941 + T10936;
  assign T10936 = {T10939, T10937};
  assign T10937 = $signed(T10938) / $signed(22'h100000);
  assign T10938 = $signed(28'h5e1d61a) * $signed(16'hffff);
  assign T10939 = T10940 ? 3'h7 : 3'h0;
  assign T10940 = T10937[6'h2b:6'h2b];
  assign T10941 = $signed(T10942) / $signed(22'h100000);
  assign T10942 = $signed(31'h3fbaa73f) * $signed(16'h0);
  assign T10943 = T10817[1'h0:1'h0];
  assign T10944 = T10817[1'h1:1'h1];
  assign T10945 = T10817[2'h2:2'h2];
  assign T10946 = T10876[6'h2e:6'h2e];
  assign T10947 = T10817[2'h3:2'h3];
  assign T10948 = {T11091, T10949};
  assign T10949 = T11090 ? T11020 : T10950;
  assign T10950 = T11019 ? T10985 : T10951;
  assign T10951 = T10984 ? T10968 : T10952;
  assign T10952 = T10967 ? twiddle4_2_17_imag : twiddle4_2_16_imag;
  assign twiddle4_2_16_imag = T10958 + T10953;
  assign T10953 = {T10956, T10954};
  assign T10954 = $signed(T10955) / $signed(22'h100000);
  assign T10955 = $signed(28'h645e9af) * $signed(16'hffff);
  assign T10956 = T10957 ? 3'h7 : 3'h0;
  assign T10957 = T10954[6'h2b:6'h2b];
  assign T10958 = $signed(T10959) / $signed(22'h100000);
  assign T10959 = $signed(31'h3fb11b47) * $signed(16'h0);
  assign twiddle4_2_17_imag = T10965 + T10960;
  assign T10960 = {T10963, T10961};
  assign T10961 = $signed(T10962) / $signed(22'h100000);
  assign T10962 = $signed(28'h6a9edc9) * $signed(16'hffff);
  assign T10963 = T10964 ? 3'h7 : 3'h0;
  assign T10964 = T10961[6'h2b:6'h2b];
  assign T10965 = $signed(T10966) / $signed(22'h100000);
  assign T10966 = $signed(31'h3fa6f228) * $signed(16'h0);
  assign T10967 = T10817[1'h0:1'h0];
  assign T10968 = T10983 ? twiddle4_2_19_imag : twiddle4_2_18_imag;
  assign twiddle4_2_18_imag = T10974 + T10969;
  assign T10969 = {T10972, T10970};
  assign T10970 = $signed(T10971) / $signed(22'h100000);
  assign T10971 = $signed(28'h70de171) * $signed(16'hffff);
  assign T10972 = T10973 ? 3'h7 : 3'h0;
  assign T10973 = T10970[6'h2b:6'h2b];
  assign T10974 = $signed(T10975) / $signed(22'h100000);
  assign T10975 = $signed(31'h3f9c2bfa) * $signed(16'h0);
  assign twiddle4_2_19_imag = T10981 + T10976;
  assign T10976 = {T10979, T10977};
  assign T10977 = $signed(T10978) / $signed(22'h100000);
  assign T10978 = $signed(28'h771c3b2) * $signed(16'hffff);
  assign T10979 = T10980 ? 3'h7 : 3'h0;
  assign T10980 = T10977[6'h2b:6'h2b];
  assign T10981 = $signed(T10982) / $signed(22'h100000);
  assign T10982 = $signed(31'h3f90c8d9) * $signed(16'h0);
  assign T10983 = T10817[1'h0:1'h0];
  assign T10984 = T10817[1'h1:1'h1];
  assign T10985 = T11018 ? T11002 : T10986;
  assign T10986 = T11001 ? twiddle4_2_21_imag : twiddle4_2_20_imag;
  assign twiddle4_2_20_imag = T10992 + T10987;
  assign T10987 = {T10990, T10988};
  assign T10988 = $signed(T10989) / $signed(22'h100000);
  assign T10989 = $signed(28'h7d59395) * $signed(16'hffff);
  assign T10990 = T10991 ? 3'h7 : 3'h0;
  assign T10991 = T10988[6'h2b:6'h2b];
  assign T10992 = $signed(T10993) / $signed(22'h100000);
  assign T10993 = $signed(31'h3f84c8e1) * $signed(16'h0);
  assign twiddle4_2_21_imag = T10999 + T10994;
  assign T10994 = {T10997, T10995};
  assign T10995 = $signed(T10996) / $signed(22'h100000);
  assign T10996 = $signed(29'h8395023) * $signed(16'hffff);
  assign T10997 = T10998 ? 2'h3 : 2'h0;
  assign T10998 = T10995[6'h2c:6'h2c];
  assign T10999 = $signed(T11000) / $signed(22'h100000);
  assign T11000 = $signed(31'h3f782c2f) * $signed(16'h0);
  assign T11001 = T10817[1'h0:1'h0];
  assign T11002 = T11017 ? twiddle4_2_23_imag : twiddle4_2_22_imag;
  assign twiddle4_2_22_imag = T11008 + T11003;
  assign T11003 = {T11006, T11004};
  assign T11004 = $signed(T11005) / $signed(22'h100000);
  assign T11005 = $signed(29'h89cf867) * $signed(16'hffff);
  assign T11006 = T11007 ? 2'h3 : 2'h0;
  assign T11007 = T11004[6'h2c:6'h2c];
  assign T11008 = $signed(T11009) / $signed(22'h100000);
  assign T11009 = $signed(31'h3f6af2e3) * $signed(16'h0);
  assign twiddle4_2_23_imag = T11015 + T11010;
  assign T11010 = {T11013, T11011};
  assign T11011 = $signed(T11012) / $signed(22'h100000);
  assign T11012 = $signed(29'h9008b6a) * $signed(16'hffff);
  assign T11013 = T11014 ? 2'h3 : 2'h0;
  assign T11014 = T11011[6'h2c:6'h2c];
  assign T11015 = $signed(T11016) / $signed(22'h100000);
  assign T11016 = $signed(31'h3f5d1d1c) * $signed(16'h0);
  assign T11017 = T10817[1'h0:1'h0];
  assign T11018 = T10817[1'h1:1'h1];
  assign T11019 = T10817[2'h2:2'h2];
  assign T11020 = T11089 ? T11055 : T11021;
  assign T11021 = T11054 ? T11038 : T11022;
  assign T11022 = T11037 ? twiddle4_2_25_imag : twiddle4_2_24_imag;
  assign twiddle4_2_24_imag = T11028 + T11023;
  assign T11023 = {T11026, T11024};
  assign T11024 = $signed(T11025) / $signed(22'h100000);
  assign T11025 = $signed(29'h9640837) * $signed(16'hffff);
  assign T11026 = T11027 ? 2'h3 : 2'h0;
  assign T11027 = T11024[6'h2c:6'h2c];
  assign T11028 = $signed(T11029) / $signed(22'h100000);
  assign T11029 = $signed(31'h3f4eaafe) * $signed(16'h0);
  assign twiddle4_2_25_imag = T11035 + T11030;
  assign T11030 = {T11033, T11031};
  assign T11031 = $signed(T11032) / $signed(22'h100000);
  assign T11032 = $signed(29'h9c76dd8) * $signed(16'hffff);
  assign T11033 = T11034 ? 2'h3 : 2'h0;
  assign T11034 = T11031[6'h2c:6'h2c];
  assign T11035 = $signed(T11036) / $signed(22'h100000);
  assign T11036 = $signed(31'h3f3f9cab) * $signed(16'h0);
  assign T11037 = T10817[1'h0:1'h0];
  assign T11038 = T11053 ? twiddle4_2_27_imag : twiddle4_2_26_imag;
  assign twiddle4_2_26_imag = T11044 + T11039;
  assign T11039 = {T11042, T11040};
  assign T11040 = $signed(T11041) / $signed(22'h100000);
  assign T11041 = $signed(29'ha2abb58) * $signed(16'hffff);
  assign T11042 = T11043 ? 2'h3 : 2'h0;
  assign T11043 = T11040[6'h2c:6'h2c];
  assign T11044 = $signed(T11045) / $signed(22'h100000);
  assign T11045 = $signed(31'h3f2ff249) * $signed(16'h0);
  assign twiddle4_2_27_imag = T11051 + T11046;
  assign T11046 = {T11049, T11047};
  assign T11047 = $signed(T11048) / $signed(22'h100000);
  assign T11048 = $signed(29'ha8defc2) * $signed(16'hffff);
  assign T11049 = T11050 ? 2'h3 : 2'h0;
  assign T11050 = T11047[6'h2c:6'h2c];
  assign T11051 = $signed(T11052) / $signed(22'h100000);
  assign T11052 = $signed(31'h3f1fabff) * $signed(16'h0);
  assign T11053 = T10817[1'h0:1'h0];
  assign T11054 = T10817[1'h1:1'h1];
  assign T11055 = T11088 ? T11072 : T11056;
  assign T11056 = T11071 ? twiddle4_2_29_imag : twiddle4_2_28_imag;
  assign twiddle4_2_28_imag = T11062 + T11057;
  assign T11057 = {T11060, T11058};
  assign T11058 = $signed(T11059) / $signed(22'h100000);
  assign T11059 = $signed(29'haf10a22) * $signed(16'hffff);
  assign T11060 = T11061 ? 2'h3 : 2'h0;
  assign T11061 = T11058[6'h2c:6'h2c];
  assign T11062 = $signed(T11063) / $signed(22'h100000);
  assign T11063 = $signed(31'h3f0ec9f4) * $signed(16'h0);
  assign twiddle4_2_29_imag = T11069 + T11064;
  assign T11064 = {T11067, T11065};
  assign T11065 = $signed(T11066) / $signed(22'h100000);
  assign T11066 = $signed(29'hb540982) * $signed(16'hffff);
  assign T11067 = T11068 ? 2'h3 : 2'h0;
  assign T11068 = T11065[6'h2c:6'h2c];
  assign T11069 = $signed(T11070) / $signed(22'h100000);
  assign T11070 = $signed(31'h3efd4c53) * $signed(16'h0);
  assign T11071 = T10817[1'h0:1'h0];
  assign T11072 = T11087 ? twiddle4_2_31_imag : twiddle4_2_30_imag;
  assign twiddle4_2_30_imag = T11078 + T11073;
  assign T11073 = {T11076, T11074};
  assign T11074 = $signed(T11075) / $signed(22'h100000);
  assign T11075 = $signed(29'hbb6ecef) * $signed(16'hffff);
  assign T11076 = T11077 ? 2'h3 : 2'h0;
  assign T11077 = T11074[6'h2c:6'h2c];
  assign T11078 = $signed(T11079) / $signed(22'h100000);
  assign T11079 = $signed(31'h3eeb3347) * $signed(16'h0);
  assign twiddle4_2_31_imag = T11085 + T11080;
  assign T11080 = {T11083, T11081};
  assign T11081 = $signed(T11082) / $signed(22'h100000);
  assign T11082 = $signed(29'hc19b374) * $signed(16'hffff);
  assign T11083 = T11084 ? 2'h3 : 2'h0;
  assign T11084 = T11081[6'h2c:6'h2c];
  assign T11085 = $signed(T11086) / $signed(22'h100000);
  assign T11086 = $signed(31'h3ed87efb) * $signed(16'h0);
  assign T11087 = T10817[1'h0:1'h0];
  assign T11088 = T10817[1'h1:1'h1];
  assign T11089 = T10817[2'h2:2'h2];
  assign T11090 = T10817[2'h3:2'h3];
  assign T11091 = T10949[6'h2e:6'h2e];
  assign T11092 = T10817[3'h4:3'h4];
  assign T11093 = {T11358, T11094};
  assign T11094 = T11357 ? T11231 : T11095;
  assign T11095 = T11230 ? T11166 : T11096;
  assign T11096 = T11165 ? T11131 : T11097;
  assign T11097 = T11130 ? T11114 : T11098;
  assign T11098 = T11113 ? twiddle4_2_33_imag : twiddle4_2_32_imag;
  assign twiddle4_2_32_imag = T11104 + T11099;
  assign T11099 = {T11102, T11100};
  assign T11100 = $signed(T11101) / $signed(22'h100000);
  assign T11101 = $signed(29'hc7c5c1e) * $signed(16'hffff);
  assign T11102 = T11103 ? 2'h3 : 2'h0;
  assign T11103 = T11100[6'h2c:6'h2c];
  assign T11104 = $signed(T11105) / $signed(22'h100000);
  assign T11105 = $signed(31'h3ec52f9f) * $signed(16'h0);
  assign twiddle4_2_33_imag = T11111 + T11106;
  assign T11106 = {T11109, T11107};
  assign T11107 = $signed(T11108) / $signed(22'h100000);
  assign T11108 = $signed(29'hcdee5f9) * $signed(16'hffff);
  assign T11109 = T11110 ? 2'h3 : 2'h0;
  assign T11110 = T11107[6'h2c:6'h2c];
  assign T11111 = $signed(T11112) / $signed(22'h100000);
  assign T11112 = $signed(31'h3eb14562) * $signed(16'h0);
  assign T11113 = T10817[1'h0:1'h0];
  assign T11114 = T11129 ? twiddle4_2_35_imag : twiddle4_2_34_imag;
  assign twiddle4_2_34_imag = T11120 + T11115;
  assign T11115 = {T11118, T11116};
  assign T11116 = $signed(T11117) / $signed(22'h100000);
  assign T11117 = $signed(29'hd415012) * $signed(16'hffff);
  assign T11118 = T11119 ? 2'h3 : 2'h0;
  assign T11119 = T11116[6'h2c:6'h2c];
  assign T11120 = $signed(T11121) / $signed(22'h100000);
  assign T11121 = $signed(31'h3e9cc076) * $signed(16'h0);
  assign twiddle4_2_35_imag = T11127 + T11122;
  assign T11122 = {T11125, T11123};
  assign T11123 = $signed(T11124) / $signed(22'h100000);
  assign T11124 = $signed(29'hda39977) * $signed(16'hffff);
  assign T11125 = T11126 ? 2'h3 : 2'h0;
  assign T11126 = T11123[6'h2c:6'h2c];
  assign T11127 = $signed(T11128) / $signed(22'h100000);
  assign T11128 = $signed(31'h3e87a10b) * $signed(16'h0);
  assign T11129 = T10817[1'h0:1'h0];
  assign T11130 = T10817[1'h1:1'h1];
  assign T11131 = T11164 ? T11148 : T11132;
  assign T11132 = T11147 ? twiddle4_2_37_imag : twiddle4_2_36_imag;
  assign twiddle4_2_36_imag = T11138 + T11133;
  assign T11133 = {T11136, T11134};
  assign T11134 = $signed(T11135) / $signed(22'h100000);
  assign T11135 = $signed(29'he05c135) * $signed(16'hffff);
  assign T11136 = T11137 ? 2'h3 : 2'h0;
  assign T11137 = T11134[6'h2c:6'h2c];
  assign T11138 = $signed(T11139) / $signed(22'h100000);
  assign T11139 = $signed(31'h3e71e758) * $signed(16'h0);
  assign twiddle4_2_37_imag = T11145 + T11140;
  assign T11140 = {T11143, T11141};
  assign T11141 = $signed(T11142) / $signed(22'h100000);
  assign T11142 = $signed(29'he67c659) * $signed(16'hffff);
  assign T11143 = T11144 ? 2'h3 : 2'h0;
  assign T11144 = T11141[6'h2c:6'h2c];
  assign T11145 = $signed(T11146) / $signed(22'h100000);
  assign T11146 = $signed(31'h3e5b9392) * $signed(16'h0);
  assign T11147 = T10817[1'h0:1'h0];
  assign T11148 = T11163 ? twiddle4_2_39_imag : twiddle4_2_38_imag;
  assign twiddle4_2_38_imag = T11154 + T11149;
  assign T11149 = {T11152, T11150};
  assign T11150 = $signed(T11151) / $signed(22'h100000);
  assign T11151 = $signed(29'hec9a7f2) * $signed(16'hffff);
  assign T11152 = T11153 ? 2'h3 : 2'h0;
  assign T11153 = T11150[6'h2c:6'h2c];
  assign T11154 = $signed(T11155) / $signed(22'h100000);
  assign T11155 = $signed(31'h3e44a5ee) * $signed(16'h0);
  assign twiddle4_2_39_imag = T11161 + T11156;
  assign T11156 = {T11159, T11157};
  assign T11157 = $signed(T11158) / $signed(22'h100000);
  assign T11158 = $signed(29'hf2b650f) * $signed(16'hffff);
  assign T11159 = T11160 ? 2'h3 : 2'h0;
  assign T11160 = T11157[6'h2c:6'h2c];
  assign T11161 = $signed(T11162) / $signed(22'h100000);
  assign T11162 = $signed(31'h3e2d1ea7) * $signed(16'h0);
  assign T11163 = T10817[1'h0:1'h0];
  assign T11164 = T10817[1'h1:1'h1];
  assign T11165 = T10817[2'h2:2'h2];
  assign T11166 = T11229 ? T11199 : T11167;
  assign T11167 = T11198 ? T11184 : T11168;
  assign T11168 = T11183 ? twiddle4_2_41_imag : twiddle4_2_40_imag;
  assign twiddle4_2_40_imag = T11174 + T11169;
  assign T11169 = {T11172, T11170};
  assign T11170 = $signed(T11171) / $signed(22'h100000);
  assign T11171 = $signed(29'hf8cfcbd) * $signed(16'hffff);
  assign T11172 = T11173 ? 2'h3 : 2'h0;
  assign T11173 = T11170[6'h2c:6'h2c];
  assign T11174 = $signed(T11175) / $signed(22'h100000);
  assign T11175 = $signed(31'h3e14fdf7) * $signed(16'h0);
  assign twiddle4_2_41_imag = T11181 + T11176;
  assign T11176 = {T11179, T11177};
  assign T11177 = $signed(T11178) / $signed(22'h100000);
  assign T11178 = $signed(29'hfee6e0d) * $signed(16'hffff);
  assign T11179 = T11180 ? 2'h3 : 2'h0;
  assign T11180 = T11177[6'h2c:6'h2c];
  assign T11181 = $signed(T11182) / $signed(22'h100000);
  assign T11182 = $signed(31'h3dfc4418) * $signed(16'h0);
  assign T11183 = T10817[1'h0:1'h0];
  assign T11184 = T11197 ? twiddle4_2_43_imag : twiddle4_2_42_imag;
  assign twiddle4_2_42_imag = T11189 + T11185;
  assign T11185 = {T11188, T11186};
  assign T11186 = $signed(T11187) / $signed(22'h100000);
  assign T11187 = $signed(30'h104fb80e) * $signed(16'hffff);
  assign T11188 = T11186[6'h2d:6'h2d];
  assign T11189 = $signed(T11190) / $signed(22'h100000);
  assign T11190 = $signed(31'h3de2f147) * $signed(16'h0);
  assign twiddle4_2_43_imag = T11195 + T11191;
  assign T11191 = {T11194, T11192};
  assign T11192 = $signed(T11193) / $signed(22'h100000);
  assign T11193 = $signed(30'h10b0d9cf) * $signed(16'hffff);
  assign T11194 = T11192[6'h2d:6'h2d];
  assign T11195 = $signed(T11196) / $signed(22'h100000);
  assign T11196 = $signed(31'h3dc905c4) * $signed(16'h0);
  assign T11197 = T10817[1'h0:1'h0];
  assign T11198 = T10817[1'h1:1'h1];
  assign T11199 = T11228 ? T11214 : T11200;
  assign T11200 = T11213 ? twiddle4_2_45_imag : twiddle4_2_44_imag;
  assign twiddle4_2_44_imag = T11205 + T11201;
  assign T11201 = {T11204, T11202};
  assign T11202 = $signed(T11203) / $signed(22'h100000);
  assign T11203 = $signed(30'h1111d262) * $signed(16'hffff);
  assign T11204 = T11202[6'h2d:6'h2d];
  assign T11205 = $signed(T11206) / $signed(22'h100000);
  assign T11206 = $signed(31'h3dae81ce) * $signed(16'h0);
  assign twiddle4_2_45_imag = T11211 + T11207;
  assign T11207 = {T11210, T11208};
  assign T11208 = $signed(T11209) / $signed(22'h100000);
  assign T11209 = $signed(30'h1172a0d7) * $signed(16'hffff);
  assign T11210 = T11208[6'h2d:6'h2d];
  assign T11211 = $signed(T11212) / $signed(22'h100000);
  assign T11212 = $signed(31'h3d9365a7) * $signed(16'h0);
  assign T11213 = T10817[1'h0:1'h0];
  assign T11214 = T11227 ? twiddle4_2_47_imag : twiddle4_2_46_imag;
  assign twiddle4_2_46_imag = T11219 + T11215;
  assign T11215 = {T11218, T11216};
  assign T11216 = $signed(T11217) / $signed(22'h100000);
  assign T11217 = $signed(30'h11d3443f) * $signed(16'hffff);
  assign T11218 = T11216[6'h2d:6'h2d];
  assign T11219 = $signed(T11220) / $signed(22'h100000);
  assign T11220 = $signed(31'h3d77b191) * $signed(16'h0);
  assign twiddle4_2_47_imag = T11225 + T11221;
  assign T11221 = {T11224, T11222};
  assign T11222 = $signed(T11223) / $signed(22'h100000);
  assign T11223 = $signed(30'h1233bbab) * $signed(16'hffff);
  assign T11224 = T11222[6'h2d:6'h2d];
  assign T11225 = $signed(T11226) / $signed(22'h100000);
  assign T11226 = $signed(31'h3d5b65d1) * $signed(16'h0);
  assign T11227 = T10817[1'h0:1'h0];
  assign T11228 = T10817[1'h1:1'h1];
  assign T11229 = T10817[2'h2:2'h2];
  assign T11230 = T10817[2'h3:2'h3];
  assign T11231 = T11356 ? T11294 : T11232;
  assign T11232 = T11293 ? T11263 : T11233;
  assign T11233 = T11262 ? T11248 : T11234;
  assign T11234 = T11247 ? twiddle4_2_49_imag : twiddle4_2_48_imag;
  assign twiddle4_2_48_imag = T11239 + T11235;
  assign T11235 = {T11238, T11236};
  assign T11236 = $signed(T11237) / $signed(22'h100000);
  assign T11237 = $signed(30'h1294062e) * $signed(16'hffff);
  assign T11238 = T11236[6'h2d:6'h2d];
  assign T11239 = $signed(T11240) / $signed(22'h100000);
  assign T11240 = $signed(31'h3d3e82ad) * $signed(16'h0);
  assign twiddle4_2_49_imag = T11245 + T11241;
  assign T11241 = {T11244, T11242};
  assign T11242 = $signed(T11243) / $signed(22'h100000);
  assign T11243 = $signed(30'h12f422da) * $signed(16'hffff);
  assign T11244 = T11242[6'h2d:6'h2d];
  assign T11245 = $signed(T11246) / $signed(22'h100000);
  assign T11246 = $signed(31'h3d21086c) * $signed(16'h0);
  assign T11247 = T10817[1'h0:1'h0];
  assign T11248 = T11261 ? twiddle4_2_51_imag : twiddle4_2_50_imag;
  assign twiddle4_2_50_imag = T11253 + T11249;
  assign T11249 = {T11252, T11250};
  assign T11250 = $signed(T11251) / $signed(22'h100000);
  assign T11251 = $signed(30'h135410c2) * $signed(16'hffff);
  assign T11252 = T11250[6'h2d:6'h2d];
  assign T11253 = $signed(T11254) / $signed(22'h100000);
  assign T11254 = $signed(31'h3d02f756) * $signed(16'h0);
  assign twiddle4_2_51_imag = T11259 + T11255;
  assign T11255 = {T11258, T11256};
  assign T11256 = $signed(T11257) / $signed(22'h100000);
  assign T11257 = $signed(30'h13b3cefa) * $signed(16'hffff);
  assign T11258 = T11256[6'h2d:6'h2d];
  assign T11259 = $signed(T11260) / $signed(22'h100000);
  assign T11260 = $signed(31'h3ce44fb6) * $signed(16'h0);
  assign T11261 = T10817[1'h0:1'h0];
  assign T11262 = T10817[1'h1:1'h1];
  assign T11263 = T11292 ? T11278 : T11264;
  assign T11264 = T11277 ? twiddle4_2_53_imag : twiddle4_2_52_imag;
  assign twiddle4_2_52_imag = T11269 + T11265;
  assign T11265 = {T11268, T11266};
  assign T11266 = $signed(T11267) / $signed(22'h100000);
  assign T11267 = $signed(30'h14135c94) * $signed(16'hffff);
  assign T11268 = T11266[6'h2d:6'h2d];
  assign T11269 = $signed(T11270) / $signed(22'h100000);
  assign T11270 = $signed(31'h3cc511d8) * $signed(16'h0);
  assign twiddle4_2_53_imag = T11275 + T11271;
  assign T11271 = {T11274, T11272};
  assign T11272 = $signed(T11273) / $signed(22'h100000);
  assign T11273 = $signed(30'h1472b8a5) * $signed(16'hffff);
  assign T11274 = T11272[6'h2d:6'h2d];
  assign T11275 = $signed(T11276) / $signed(22'h100000);
  assign T11276 = $signed(31'h3ca53e08) * $signed(16'h0);
  assign T11277 = T10817[1'h0:1'h0];
  assign T11278 = T11291 ? twiddle4_2_55_imag : twiddle4_2_54_imag;
  assign twiddle4_2_54_imag = T11283 + T11279;
  assign T11279 = {T11282, T11280};
  assign T11280 = $signed(T11281) / $signed(22'h100000);
  assign T11281 = $signed(30'h14d1e242) * $signed(16'hffff);
  assign T11282 = T11280[6'h2d:6'h2d];
  assign T11283 = $signed(T11284) / $signed(22'h100000);
  assign T11284 = $signed(31'h3c84d496) * $signed(16'h0);
  assign twiddle4_2_55_imag = T11289 + T11285;
  assign T11285 = {T11288, T11286};
  assign T11286 = $signed(T11287) / $signed(22'h100000);
  assign T11287 = $signed(30'h1530d880) * $signed(16'hffff);
  assign T11288 = T11286[6'h2d:6'h2d];
  assign T11289 = $signed(T11290) / $signed(22'h100000);
  assign T11290 = $signed(31'h3c63d5d0) * $signed(16'h0);
  assign T11291 = T10817[1'h0:1'h0];
  assign T11292 = T10817[1'h1:1'h1];
  assign T11293 = T10817[2'h2:2'h2];
  assign T11294 = T11355 ? T11325 : T11295;
  assign T11295 = T11324 ? T11310 : T11296;
  assign T11296 = T11309 ? twiddle4_2_57_imag : twiddle4_2_56_imag;
  assign twiddle4_2_56_imag = T11301 + T11297;
  assign T11297 = {T11300, T11298};
  assign T11298 = $signed(T11299) / $signed(22'h100000);
  assign T11299 = $signed(30'h158f9a75) * $signed(16'hffff);
  assign T11300 = T11298[6'h2d:6'h2d];
  assign T11301 = $signed(T11302) / $signed(22'h100000);
  assign T11302 = $signed(31'h3c424209) * $signed(16'h0);
  assign twiddle4_2_57_imag = T11307 + T11303;
  assign T11303 = {T11306, T11304};
  assign T11304 = $signed(T11305) / $signed(22'h100000);
  assign T11305 = $signed(30'h15ee2737) * $signed(16'hffff);
  assign T11306 = T11304[6'h2d:6'h2d];
  assign T11307 = $signed(T11308) / $signed(22'h100000);
  assign T11308 = $signed(31'h3c201994) * $signed(16'h0);
  assign T11309 = T10817[1'h0:1'h0];
  assign T11310 = T11323 ? twiddle4_2_59_imag : twiddle4_2_58_imag;
  assign twiddle4_2_58_imag = T11315 + T11311;
  assign T11311 = {T11314, T11312};
  assign T11312 = $signed(T11313) / $signed(22'h100000);
  assign T11313 = $signed(30'h164c7ddd) * $signed(16'hffff);
  assign T11314 = T11312[6'h2d:6'h2d];
  assign T11315 = $signed(T11316) / $signed(22'h100000);
  assign T11316 = $signed(31'h3bfd5cc4) * $signed(16'h0);
  assign twiddle4_2_59_imag = T11321 + T11317;
  assign T11317 = {T11320, T11318};
  assign T11318 = $signed(T11319) / $signed(22'h100000);
  assign T11319 = $signed(30'h16aa9d7d) * $signed(16'hffff);
  assign T11320 = T11318[6'h2d:6'h2d];
  assign T11321 = $signed(T11322) / $signed(22'h100000);
  assign T11322 = $signed(31'h3bda0bef) * $signed(16'h0);
  assign T11323 = T10817[1'h0:1'h0];
  assign T11324 = T10817[1'h1:1'h1];
  assign T11325 = T11354 ? T11340 : T11326;
  assign T11326 = T11339 ? twiddle4_2_61_imag : twiddle4_2_60_imag;
  assign twiddle4_2_60_imag = T11331 + T11327;
  assign T11327 = {T11330, T11328};
  assign T11328 = $signed(T11329) / $signed(22'h100000);
  assign T11329 = $signed(30'h17088530) * $signed(16'hffff);
  assign T11330 = T11328[6'h2d:6'h2d];
  assign T11331 = $signed(T11332) / $signed(22'h100000);
  assign T11332 = $signed(31'h3bb6276d) * $signed(16'h0);
  assign twiddle4_2_61_imag = T11337 + T11333;
  assign T11333 = {T11336, T11334};
  assign T11334 = $signed(T11335) / $signed(22'h100000);
  assign T11335 = $signed(30'h1766340f) * $signed(16'hffff);
  assign T11336 = T11334[6'h2d:6'h2d];
  assign T11337 = $signed(T11338) / $signed(22'h100000);
  assign T11338 = $signed(31'h3b91af96) * $signed(16'h0);
  assign T11339 = T10817[1'h0:1'h0];
  assign T11340 = T11353 ? twiddle4_2_63_imag : twiddle4_2_62_imag;
  assign twiddle4_2_62_imag = T11345 + T11341;
  assign T11341 = {T11344, T11342};
  assign T11342 = $signed(T11343) / $signed(22'h100000);
  assign T11343 = $signed(30'h17c3a931) * $signed(16'hffff);
  assign T11344 = T11342[6'h2d:6'h2d];
  assign T11345 = $signed(T11346) / $signed(22'h100000);
  assign T11346 = $signed(31'h3b6ca4c4) * $signed(16'h0);
  assign twiddle4_2_63_imag = T11351 + T11347;
  assign T11347 = {T11350, T11348};
  assign T11348 = $signed(T11349) / $signed(22'h100000);
  assign T11349 = $signed(30'h1820e3b0) * $signed(16'hffff);
  assign T11350 = T11348[6'h2d:6'h2d];
  assign T11351 = $signed(T11352) / $signed(22'h100000);
  assign T11352 = $signed(31'h3b470752) * $signed(16'h0);
  assign T11353 = T10817[1'h0:1'h0];
  assign T11354 = T10817[1'h1:1'h1];
  assign T11355 = T10817[2'h2:2'h2];
  assign T11356 = T10817[2'h3:2'h3];
  assign T11357 = T10817[3'h4:3'h4];
  assign T11358 = T11094[6'h2e:6'h2e];
  assign T11359 = T10817[3'h5:3'h5];
  assign T11360 = {T11787, T11361};
  assign T11361 = T11786 ? T11596 : T11362;
  assign T11362 = T11595 ? T11489 : T11363;
  assign T11363 = T11488 ? T11426 : T11364;
  assign T11364 = T11425 ? T11395 : T11365;
  assign T11365 = T11394 ? T11380 : T11366;
  assign T11366 = T11379 ? twiddle4_2_65_imag : twiddle4_2_64_imag;
  assign twiddle4_2_64_imag = T11371 + T11367;
  assign T11367 = {T11370, T11368};
  assign T11368 = $signed(T11369) / $signed(22'h100000);
  assign T11369 = $signed(30'h187de2a6) * $signed(16'hffff);
  assign T11370 = T11368[6'h2d:6'h2d];
  assign T11371 = $signed(T11372) / $signed(22'h100000);
  assign T11372 = $signed(31'h3b20d79e) * $signed(16'h0);
  assign twiddle4_2_65_imag = T11377 + T11373;
  assign T11373 = {T11376, T11374};
  assign T11374 = $signed(T11375) / $signed(22'h100000);
  assign T11375 = $signed(30'h18daa52e) * $signed(16'hffff);
  assign T11376 = T11374[6'h2d:6'h2d];
  assign T11377 = $signed(T11378) / $signed(22'h100000);
  assign T11378 = $signed(31'h3afa1605) * $signed(16'h0);
  assign T11379 = T10817[1'h0:1'h0];
  assign T11380 = T11393 ? twiddle4_2_67_imag : twiddle4_2_66_imag;
  assign twiddle4_2_66_imag = T11385 + T11381;
  assign T11381 = {T11384, T11382};
  assign T11382 = $signed(T11383) / $signed(22'h100000);
  assign T11383 = $signed(30'h19372a63) * $signed(16'hffff);
  assign T11384 = T11382[6'h2d:6'h2d];
  assign T11385 = $signed(T11386) / $signed(22'h100000);
  assign T11386 = $signed(31'h3ad2c2e7) * $signed(16'h0);
  assign twiddle4_2_67_imag = T11391 + T11387;
  assign T11387 = {T11390, T11388};
  assign T11388 = $signed(T11389) / $signed(22'h100000);
  assign T11389 = $signed(30'h19937161) * $signed(16'hffff);
  assign T11390 = T11388[6'h2d:6'h2d];
  assign T11391 = $signed(T11392) / $signed(22'h100000);
  assign T11392 = $signed(31'h3aaadea5) * $signed(16'h0);
  assign T11393 = T10817[1'h0:1'h0];
  assign T11394 = T10817[1'h1:1'h1];
  assign T11395 = T11424 ? T11410 : T11396;
  assign T11396 = T11409 ? twiddle4_2_69_imag : twiddle4_2_68_imag;
  assign twiddle4_2_68_imag = T11401 + T11397;
  assign T11397 = {T11400, T11398};
  assign T11398 = $signed(T11399) / $signed(22'h100000);
  assign T11399 = $signed(30'h19ef7943) * $signed(16'hffff);
  assign T11400 = T11398[6'h2d:6'h2d];
  assign T11401 = $signed(T11402) / $signed(22'h100000);
  assign T11402 = $signed(31'h3a8269a2) * $signed(16'h0);
  assign twiddle4_2_69_imag = T11407 + T11403;
  assign T11403 = {T11406, T11404};
  assign T11404 = $signed(T11405) / $signed(22'h100000);
  assign T11405 = $signed(30'h1a4b4127) * $signed(16'hffff);
  assign T11406 = T11404[6'h2d:6'h2d];
  assign T11407 = $signed(T11408) / $signed(22'h100000);
  assign T11408 = $signed(31'h3a596441) * $signed(16'h0);
  assign T11409 = T10817[1'h0:1'h0];
  assign T11410 = T11423 ? twiddle4_2_71_imag : twiddle4_2_70_imag;
  assign twiddle4_2_70_imag = T11415 + T11411;
  assign T11411 = {T11414, T11412};
  assign T11412 = $signed(T11413) / $signed(22'h100000);
  assign T11413 = $signed(30'h1aa6c82b) * $signed(16'hffff);
  assign T11414 = T11412[6'h2d:6'h2d];
  assign T11415 = $signed(T11416) / $signed(22'h100000);
  assign T11416 = $signed(31'h3a2fcee8) * $signed(16'h0);
  assign twiddle4_2_71_imag = T11421 + T11417;
  assign T11417 = {T11420, T11418};
  assign T11418 = $signed(T11419) / $signed(22'h100000);
  assign T11419 = $signed(30'h1b020d6c) * $signed(16'hffff);
  assign T11420 = T11418[6'h2d:6'h2d];
  assign T11421 = $signed(T11422) / $signed(22'h100000);
  assign T11422 = $signed(31'h3a05a9fd) * $signed(16'h0);
  assign T11423 = T10817[1'h0:1'h0];
  assign T11424 = T10817[1'h1:1'h1];
  assign T11425 = T10817[2'h2:2'h2];
  assign T11426 = T11487 ? T11457 : T11427;
  assign T11427 = T11456 ? T11442 : T11428;
  assign T11428 = T11441 ? twiddle4_2_73_imag : twiddle4_2_72_imag;
  assign twiddle4_2_72_imag = T11433 + T11429;
  assign T11429 = {T11432, T11430};
  assign T11430 = $signed(T11431) / $signed(22'h100000);
  assign T11431 = $signed(30'h1b5d1009) * $signed(16'hffff);
  assign T11432 = T11430[6'h2d:6'h2d];
  assign T11433 = $signed(T11434) / $signed(22'h100000);
  assign T11434 = $signed(31'h39daf5e8) * $signed(16'h0);
  assign twiddle4_2_73_imag = T11439 + T11435;
  assign T11435 = {T11438, T11436};
  assign T11436 = $signed(T11437) / $signed(22'h100000);
  assign T11437 = $signed(30'h1bb7cf23) * $signed(16'hffff);
  assign T11438 = T11436[6'h2d:6'h2d];
  assign T11439 = $signed(T11440) / $signed(22'h100000);
  assign T11440 = $signed(31'h39afb313) * $signed(16'h0);
  assign T11441 = T10817[1'h0:1'h0];
  assign T11442 = T11455 ? twiddle4_2_75_imag : twiddle4_2_74_imag;
  assign twiddle4_2_74_imag = T11447 + T11443;
  assign T11443 = {T11446, T11444};
  assign T11444 = $signed(T11445) / $signed(22'h100000);
  assign T11445 = $signed(30'h1c1249d8) * $signed(16'hffff);
  assign T11446 = T11444[6'h2d:6'h2d];
  assign T11447 = $signed(T11448) / $signed(22'h100000);
  assign T11448 = $signed(31'h3983e1e7) * $signed(16'h0);
  assign twiddle4_2_75_imag = T11453 + T11449;
  assign T11449 = {T11452, T11450};
  assign T11450 = $signed(T11451) / $signed(22'h100000);
  assign T11451 = $signed(30'h1c6c7f49) * $signed(16'hffff);
  assign T11452 = T11450[6'h2d:6'h2d];
  assign T11453 = $signed(T11454) / $signed(22'h100000);
  assign T11454 = $signed(31'h395782d3) * $signed(16'h0);
  assign T11455 = T10817[1'h0:1'h0];
  assign T11456 = T10817[1'h1:1'h1];
  assign T11457 = T11486 ? T11472 : T11458;
  assign T11458 = T11471 ? twiddle4_2_77_imag : twiddle4_2_76_imag;
  assign twiddle4_2_76_imag = T11463 + T11459;
  assign T11459 = {T11462, T11460};
  assign T11460 = $signed(T11461) / $signed(22'h100000);
  assign T11461 = $signed(30'h1cc66e99) * $signed(16'hffff);
  assign T11462 = T11460[6'h2d:6'h2d];
  assign T11463 = $signed(T11464) / $signed(22'h100000);
  assign T11464 = $signed(31'h392a9642) * $signed(16'h0);
  assign twiddle4_2_77_imag = T11469 + T11465;
  assign T11465 = {T11468, T11466};
  assign T11466 = $signed(T11467) / $signed(22'h100000);
  assign T11467 = $signed(30'h1d2016e8) * $signed(16'hffff);
  assign T11468 = T11466[6'h2d:6'h2d];
  assign T11469 = $signed(T11470) / $signed(22'h100000);
  assign T11470 = $signed(31'h38fd1ca4) * $signed(16'h0);
  assign T11471 = T10817[1'h0:1'h0];
  assign T11472 = T11485 ? twiddle4_2_79_imag : twiddle4_2_78_imag;
  assign twiddle4_2_78_imag = T11477 + T11473;
  assign T11473 = {T11476, T11474};
  assign T11474 = $signed(T11475) / $signed(22'h100000);
  assign T11475 = $signed(30'h1d79775b) * $signed(16'hffff);
  assign T11476 = T11474[6'h2d:6'h2d];
  assign T11477 = $signed(T11478) / $signed(22'h100000);
  assign T11478 = $signed(31'h38cf1669) * $signed(16'h0);
  assign twiddle4_2_79_imag = T11483 + T11479;
  assign T11479 = {T11482, T11480};
  assign T11480 = $signed(T11481) / $signed(22'h100000);
  assign T11481 = $signed(30'h1dd28f14) * $signed(16'hffff);
  assign T11482 = T11480[6'h2d:6'h2d];
  assign T11483 = $signed(T11484) / $signed(22'h100000);
  assign T11484 = $signed(31'h38a08402) * $signed(16'h0);
  assign T11485 = T10817[1'h0:1'h0];
  assign T11486 = T10817[1'h1:1'h1];
  assign T11487 = T10817[2'h2:2'h2];
  assign T11488 = T10817[2'h3:2'h3];
  assign T11489 = T11594 ? T11548 : T11490;
  assign T11490 = T11547 ? T11521 : T11491;
  assign T11491 = T11520 ? T11506 : T11492;
  assign T11492 = T11505 ? twiddle4_2_81_imag : twiddle4_2_80_imag;
  assign twiddle4_2_80_imag = T11497 + T11493;
  assign T11493 = {T11496, T11494};
  assign T11494 = $signed(T11495) / $signed(22'h100000);
  assign T11495 = $signed(30'h1e2b5d38) * $signed(16'hffff);
  assign T11496 = T11494[6'h2d:6'h2d];
  assign T11497 = $signed(T11498) / $signed(22'h100000);
  assign T11498 = $signed(31'h387165e3) * $signed(16'h0);
  assign twiddle4_2_81_imag = T11503 + T11499;
  assign T11499 = {T11502, T11500};
  assign T11500 = $signed(T11501) / $signed(22'h100000);
  assign T11501 = $signed(30'h1e83e0ea) * $signed(16'hffff);
  assign T11502 = T11500[6'h2d:6'h2d];
  assign T11503 = $signed(T11504) / $signed(22'h100000);
  assign T11504 = $signed(31'h3841bc7f) * $signed(16'h0);
  assign T11505 = T10817[1'h0:1'h0];
  assign T11506 = T11519 ? twiddle4_2_83_imag : twiddle4_2_82_imag;
  assign twiddle4_2_82_imag = T11511 + T11507;
  assign T11507 = {T11510, T11508};
  assign T11508 = $signed(T11509) / $signed(22'h100000);
  assign T11509 = $signed(30'h1edc1952) * $signed(16'hffff);
  assign T11510 = T11508[6'h2d:6'h2d];
  assign T11511 = $signed(T11512) / $signed(22'h100000);
  assign T11512 = $signed(31'h3811884c) * $signed(16'h0);
  assign twiddle4_2_83_imag = T11517 + T11513;
  assign T11513 = {T11516, T11514};
  assign T11514 = $signed(T11515) / $signed(22'h100000);
  assign T11515 = $signed(30'h1f340596) * $signed(16'hffff);
  assign T11516 = T11514[6'h2d:6'h2d];
  assign T11517 = $signed(T11518) / $signed(22'h100000);
  assign T11518 = $signed(31'h37e0c9c2) * $signed(16'h0);
  assign T11519 = T10817[1'h0:1'h0];
  assign T11520 = T10817[1'h1:1'h1];
  assign T11521 = T11546 ? T11536 : T11522;
  assign T11522 = T11535 ? twiddle4_2_85_imag : twiddle4_2_84_imag;
  assign twiddle4_2_84_imag = T11527 + T11523;
  assign T11523 = {T11526, T11524};
  assign T11524 = $signed(T11525) / $signed(22'h100000);
  assign T11525 = $signed(30'h1f8ba4db) * $signed(16'hffff);
  assign T11526 = T11524[6'h2d:6'h2d];
  assign T11527 = $signed(T11528) / $signed(22'h100000);
  assign T11528 = $signed(31'h37af8158) * $signed(16'h0);
  assign twiddle4_2_85_imag = T11533 + T11529;
  assign T11529 = {T11532, T11530};
  assign T11530 = $signed(T11531) / $signed(22'h100000);
  assign T11531 = $signed(30'h1fe2f64b) * $signed(16'hffff);
  assign T11532 = T11530[6'h2d:6'h2d];
  assign T11533 = $signed(T11534) / $signed(22'h100000);
  assign T11534 = $signed(31'h377daf89) * $signed(16'h0);
  assign T11535 = T10817[1'h0:1'h0];
  assign T11536 = T11545 ? twiddle4_2_87_imag : twiddle4_2_86_imag;
  assign twiddle4_2_86_imag = T11539 + T11537;
  assign T11537 = $signed(T11538) / $signed(22'h100000);
  assign T11538 = $signed(31'h2039f90e) * $signed(16'hffff);
  assign T11539 = $signed(T11540) / $signed(22'h100000);
  assign T11540 = $signed(31'h374b54ce) * $signed(16'h0);
  assign twiddle4_2_87_imag = T11543 + T11541;
  assign T11541 = $signed(T11542) / $signed(22'h100000);
  assign T11542 = $signed(31'h2090ac4d) * $signed(16'hffff);
  assign T11543 = $signed(T11544) / $signed(22'h100000);
  assign T11544 = $signed(31'h371871a4) * $signed(16'h0);
  assign T11545 = T10817[1'h0:1'h0];
  assign T11546 = T10817[1'h1:1'h1];
  assign T11547 = T10817[2'h2:2'h2];
  assign T11548 = T11593 ? T11571 : T11549;
  assign T11549 = T11570 ? T11560 : T11550;
  assign T11550 = T11559 ? twiddle4_2_89_imag : twiddle4_2_88_imag;
  assign twiddle4_2_88_imag = T11553 + T11551;
  assign T11551 = $signed(T11552) / $signed(22'h100000);
  assign T11552 = $signed(31'h20e70f32) * $signed(16'hffff);
  assign T11553 = $signed(T11554) / $signed(22'h100000);
  assign T11554 = $signed(31'h36e5068a) * $signed(16'h0);
  assign twiddle4_2_89_imag = T11557 + T11555;
  assign T11555 = $signed(T11556) / $signed(22'h100000);
  assign T11556 = $signed(31'h213d20e8) * $signed(16'hffff);
  assign T11557 = $signed(T11558) / $signed(22'h100000);
  assign T11558 = $signed(31'h36b113fd) * $signed(16'h0);
  assign T11559 = T10817[1'h0:1'h0];
  assign T11560 = T11569 ? twiddle4_2_91_imag : twiddle4_2_90_imag;
  assign twiddle4_2_90_imag = T11563 + T11561;
  assign T11561 = $signed(T11562) / $signed(22'h100000);
  assign T11562 = $signed(31'h2192e09a) * $signed(16'hffff);
  assign T11563 = $signed(T11564) / $signed(22'h100000);
  assign T11564 = $signed(31'h367c9a7d) * $signed(16'h0);
  assign twiddle4_2_91_imag = T11567 + T11565;
  assign T11565 = $signed(T11566) / $signed(22'h100000);
  assign T11566 = $signed(31'h21e84d76) * $signed(16'hffff);
  assign T11567 = $signed(T11568) / $signed(22'h100000);
  assign T11568 = $signed(31'h36479a8e) * $signed(16'h0);
  assign T11569 = T10817[1'h0:1'h0];
  assign T11570 = T10817[1'h1:1'h1];
  assign T11571 = T11592 ? T11582 : T11572;
  assign T11572 = T11581 ? twiddle4_2_93_imag : twiddle4_2_92_imag;
  assign twiddle4_2_92_imag = T11575 + T11573;
  assign T11573 = $signed(T11574) / $signed(22'h100000);
  assign T11574 = $signed(31'h223d66a8) * $signed(16'hffff);
  assign T11575 = $signed(T11576) / $signed(22'h100000);
  assign T11576 = $signed(31'h361214b0) * $signed(16'h0);
  assign twiddle4_2_93_imag = T11579 + T11577;
  assign T11577 = $signed(T11578) / $signed(22'h100000);
  assign T11578 = $signed(31'h22922b5e) * $signed(16'hffff);
  assign T11579 = $signed(T11580) / $signed(22'h100000);
  assign T11580 = $signed(31'h35dc0968) * $signed(16'h0);
  assign T11581 = T10817[1'h0:1'h0];
  assign T11582 = T11591 ? twiddle4_2_95_imag : twiddle4_2_94_imag;
  assign twiddle4_2_94_imag = T11585 + T11583;
  assign T11583 = $signed(T11584) / $signed(22'h100000);
  assign T11584 = $signed(31'h22e69ac7) * $signed(16'hffff);
  assign T11585 = $signed(T11586) / $signed(22'h100000);
  assign T11586 = $signed(31'h35a5793c) * $signed(16'h0);
  assign twiddle4_2_95_imag = T11589 + T11587;
  assign T11587 = $signed(T11588) / $signed(22'h100000);
  assign T11588 = $signed(31'h233ab413) * $signed(16'hffff);
  assign T11589 = $signed(T11590) / $signed(22'h100000);
  assign T11590 = $signed(31'h356e64b2) * $signed(16'h0);
  assign T11591 = T10817[1'h0:1'h0];
  assign T11592 = T10817[1'h1:1'h1];
  assign T11593 = T10817[2'h2:2'h2];
  assign T11594 = T10817[2'h3:2'h3];
  assign T11595 = T10817[3'h4:3'h4];
  assign T11596 = T11785 ? T11691 : T11597;
  assign T11597 = T11690 ? T11644 : T11598;
  assign T11598 = T11643 ? T11621 : T11599;
  assign T11599 = T11620 ? T11610 : T11600;
  assign T11600 = T11609 ? twiddle4_2_97_imag : twiddle4_2_96_imag;
  assign twiddle4_2_96_imag = T11603 + T11601;
  assign T11601 = $signed(T11602) / $signed(22'h100000);
  assign T11602 = $signed(31'h238e7673) * $signed(16'hffff);
  assign T11603 = $signed(T11604) / $signed(22'h100000);
  assign T11604 = $signed(31'h3536cc52) * $signed(16'h0);
  assign twiddle4_2_97_imag = T11607 + T11605;
  assign T11605 = $signed(T11606) / $signed(22'h100000);
  assign T11606 = $signed(31'h23e1e117) * $signed(16'hffff);
  assign T11607 = $signed(T11608) / $signed(22'h100000);
  assign T11608 = $signed(31'h34feb0a5) * $signed(16'h0);
  assign T11609 = T10817[1'h0:1'h0];
  assign T11610 = T11619 ? twiddle4_2_99_imag : twiddle4_2_98_imag;
  assign twiddle4_2_98_imag = T11613 + T11611;
  assign T11611 = $signed(T11612) / $signed(22'h100000);
  assign T11612 = $signed(31'h2434f332) * $signed(16'hffff);
  assign T11613 = $signed(T11614) / $signed(22'h100000);
  assign T11614 = $signed(31'h34c61236) * $signed(16'h0);
  assign twiddle4_2_99_imag = T11617 + T11615;
  assign T11615 = $signed(T11616) / $signed(22'h100000);
  assign T11616 = $signed(31'h2487abf7) * $signed(16'hffff);
  assign T11617 = $signed(T11618) / $signed(22'h100000);
  assign T11618 = $signed(31'h348cf190) * $signed(16'h0);
  assign T11619 = T10817[1'h0:1'h0];
  assign T11620 = T10817[1'h1:1'h1];
  assign T11621 = T11642 ? T11632 : T11622;
  assign T11622 = T11631 ? twiddle4_2_101_imag : twiddle4_2_100_imag;
  assign twiddle4_2_100_imag = T11625 + T11623;
  assign T11623 = $signed(T11624) / $signed(22'h100000);
  assign T11624 = $signed(31'h24da0a99) * $signed(16'hffff);
  assign T11625 = $signed(T11626) / $signed(22'h100000);
  assign T11626 = $signed(31'h34534f40) * $signed(16'h0);
  assign twiddle4_2_101_imag = T11629 + T11627;
  assign T11627 = $signed(T11628) / $signed(22'h100000);
  assign T11628 = $signed(31'h252c0e4e) * $signed(16'hffff);
  assign T11629 = $signed(T11630) / $signed(22'h100000);
  assign T11630 = $signed(31'h34192bd5) * $signed(16'h0);
  assign T11631 = T10817[1'h0:1'h0];
  assign T11632 = T11641 ? twiddle4_2_103_imag : twiddle4_2_102_imag;
  assign twiddle4_2_102_imag = T11635 + T11633;
  assign T11633 = $signed(T11634) / $signed(22'h100000);
  assign T11634 = $signed(31'h257db64b) * $signed(16'hffff);
  assign T11635 = $signed(T11636) / $signed(22'h100000);
  assign T11636 = $signed(31'h33de87de) * $signed(16'h0);
  assign twiddle4_2_103_imag = T11639 + T11637;
  assign T11637 = $signed(T11638) / $signed(22'h100000);
  assign T11638 = $signed(31'h25cf01c7) * $signed(16'hffff);
  assign T11639 = $signed(T11640) / $signed(22'h100000);
  assign T11640 = $signed(31'h33a363eb) * $signed(16'h0);
  assign T11641 = T10817[1'h0:1'h0];
  assign T11642 = T10817[1'h1:1'h1];
  assign T11643 = T10817[2'h2:2'h2];
  assign T11644 = T11689 ? T11667 : T11645;
  assign T11645 = T11666 ? T11656 : T11646;
  assign T11646 = T11655 ? twiddle4_2_105_imag : twiddle4_2_104_imag;
  assign twiddle4_2_104_imag = T11649 + T11647;
  assign T11647 = $signed(T11648) / $signed(22'h100000);
  assign T11648 = $signed(31'h261feff9) * $signed(16'hffff);
  assign T11649 = $signed(T11650) / $signed(22'h100000);
  assign T11650 = $signed(31'h3367c08f) * $signed(16'h0);
  assign twiddle4_2_105_imag = T11653 + T11651;
  assign T11651 = $signed(T11652) / $signed(22'h100000);
  assign T11652 = $signed(31'h2670801a) * $signed(16'hffff);
  assign T11653 = $signed(T11654) / $signed(22'h100000);
  assign T11654 = $signed(31'h332b9e5d) * $signed(16'h0);
  assign T11655 = T10817[1'h0:1'h0];
  assign T11656 = T11665 ? twiddle4_2_107_imag : twiddle4_2_106_imag;
  assign twiddle4_2_106_imag = T11659 + T11657;
  assign T11657 = $signed(T11658) / $signed(22'h100000);
  assign T11658 = $signed(31'h26c0b162) * $signed(16'hffff);
  assign T11659 = $signed(T11660) / $signed(22'h100000);
  assign T11660 = $signed(31'h32eefde9) * $signed(16'h0);
  assign twiddle4_2_107_imag = T11663 + T11661;
  assign T11661 = $signed(T11662) / $signed(22'h100000);
  assign T11662 = $signed(31'h2710830b) * $signed(16'hffff);
  assign T11663 = $signed(T11664) / $signed(22'h100000);
  assign T11664 = $signed(31'h32b1dfc9) * $signed(16'h0);
  assign T11665 = T10817[1'h0:1'h0];
  assign T11666 = T10817[1'h1:1'h1];
  assign T11667 = T11688 ? T11678 : T11668;
  assign T11668 = T11677 ? twiddle4_2_109_imag : twiddle4_2_108_imag;
  assign twiddle4_2_108_imag = T11671 + T11669;
  assign T11669 = $signed(T11670) / $signed(22'h100000);
  assign T11670 = $signed(31'h275ff452) * $signed(16'hffff);
  assign T11671 = $signed(T11672) / $signed(22'h100000);
  assign T11672 = $signed(31'h32744493) * $signed(16'h0);
  assign twiddle4_2_109_imag = T11675 + T11673;
  assign T11673 = $signed(T11674) / $signed(22'h100000);
  assign T11674 = $signed(31'h27af0471) * $signed(16'hffff);
  assign T11675 = $signed(T11676) / $signed(22'h100000);
  assign T11676 = $signed(31'h32362cdf) * $signed(16'h0);
  assign T11677 = T10817[1'h0:1'h0];
  assign T11678 = T11687 ? twiddle4_2_111_imag : twiddle4_2_110_imag;
  assign twiddle4_2_110_imag = T11681 + T11679;
  assign T11679 = $signed(T11680) / $signed(22'h100000);
  assign T11680 = $signed(31'h27fdb2a6) * $signed(16'hffff);
  assign T11681 = $signed(T11682) / $signed(22'h100000);
  assign T11682 = $signed(31'h31f79947) * $signed(16'h0);
  assign twiddle4_2_111_imag = T11685 + T11683;
  assign T11683 = $signed(T11684) / $signed(22'h100000);
  assign T11684 = $signed(31'h284bfe2f) * $signed(16'hffff);
  assign T11685 = $signed(T11686) / $signed(22'h100000);
  assign T11686 = $signed(31'h31b88a66) * $signed(16'h0);
  assign T11687 = T10817[1'h0:1'h0];
  assign T11688 = T10817[1'h1:1'h1];
  assign T11689 = T10817[2'h2:2'h2];
  assign T11690 = T10817[2'h3:2'h3];
  assign T11691 = T11784 ? T11738 : T11692;
  assign T11692 = T11737 ? T11715 : T11693;
  assign T11693 = T11714 ? T11704 : T11694;
  assign T11694 = T11703 ? twiddle4_2_113_imag : twiddle4_2_112_imag;
  assign twiddle4_2_112_imag = T11697 + T11695;
  assign T11695 = $signed(T11696) / $signed(22'h100000);
  assign T11696 = $signed(31'h2899e64a) * $signed(16'hffff);
  assign T11697 = $signed(T11698) / $signed(22'h100000);
  assign T11698 = $signed(31'h317900d6) * $signed(16'h0);
  assign twiddle4_2_113_imag = T11701 + T11699;
  assign T11699 = $signed(T11700) / $signed(22'h100000);
  assign T11700 = $signed(31'h28e76a37) * $signed(16'hffff);
  assign T11701 = $signed(T11702) / $signed(22'h100000);
  assign T11702 = $signed(31'h3138fd34) * $signed(16'h0);
  assign T11703 = T10817[1'h0:1'h0];
  assign T11704 = T11713 ? twiddle4_2_115_imag : twiddle4_2_114_imag;
  assign twiddle4_2_114_imag = T11707 + T11705;
  assign T11705 = $signed(T11706) / $signed(22'h100000);
  assign T11706 = $signed(31'h29348937) * $signed(16'hffff);
  assign T11707 = $signed(T11708) / $signed(22'h100000);
  assign T11708 = $signed(31'h30f8801f) * $signed(16'h0);
  assign twiddle4_2_115_imag = T11711 + T11709;
  assign T11709 = $signed(T11710) / $signed(22'h100000);
  assign T11710 = $signed(31'h2981428b) * $signed(16'hffff);
  assign T11711 = $signed(T11712) / $signed(22'h100000);
  assign T11712 = $signed(31'h30b78a35) * $signed(16'h0);
  assign T11713 = T10817[1'h0:1'h0];
  assign T11714 = T10817[1'h1:1'h1];
  assign T11715 = T11736 ? T11726 : T11716;
  assign T11716 = T11725 ? twiddle4_2_117_imag : twiddle4_2_116_imag;
  assign twiddle4_2_116_imag = T11719 + T11717;
  assign T11717 = $signed(T11718) / $signed(22'h100000);
  assign T11718 = $signed(31'h29cd9577) * $signed(16'hffff);
  assign T11719 = $signed(T11720) / $signed(22'h100000);
  assign T11720 = $signed(31'h30761c17) * $signed(16'h0);
  assign twiddle4_2_117_imag = T11723 + T11721;
  assign T11721 = $signed(T11722) / $signed(22'h100000);
  assign T11722 = $signed(31'h2a19813e) * $signed(16'hffff);
  assign T11723 = $signed(T11724) / $signed(22'h100000);
  assign T11724 = $signed(31'h30343667) * $signed(16'h0);
  assign T11725 = T10817[1'h0:1'h0];
  assign T11726 = T11735 ? twiddle4_2_119_imag : twiddle4_2_118_imag;
  assign twiddle4_2_118_imag = T11729 + T11727;
  assign T11727 = $signed(T11728) / $signed(22'h100000);
  assign T11728 = $signed(31'h2a650525) * $signed(16'hffff);
  assign T11729 = $signed(T11730) / $signed(22'h100000);
  assign T11730 = $signed(31'h2ff1d9c6) * $signed(16'h0);
  assign twiddle4_2_119_imag = T11733 + T11731;
  assign T11731 = $signed(T11732) / $signed(22'h100000);
  assign T11732 = $signed(31'h2ab02071) * $signed(16'hffff);
  assign T11733 = $signed(T11734) / $signed(22'h100000);
  assign T11734 = $signed(31'h2faf06d9) * $signed(16'h0);
  assign T11735 = T10817[1'h0:1'h0];
  assign T11736 = T10817[1'h1:1'h1];
  assign T11737 = T10817[2'h2:2'h2];
  assign T11738 = T11783 ? T11761 : T11739;
  assign T11739 = T11760 ? T11750 : T11740;
  assign T11740 = T11749 ? twiddle4_2_121_imag : twiddle4_2_120_imag;
  assign twiddle4_2_120_imag = T11743 + T11741;
  assign T11741 = $signed(T11742) / $signed(22'h100000);
  assign T11742 = $signed(31'h2afad269) * $signed(16'hffff);
  assign T11743 = $signed(T11744) / $signed(22'h100000);
  assign T11744 = $signed(31'h2f6bbe44) * $signed(16'h0);
  assign twiddle4_2_121_imag = T11747 + T11745;
  assign T11745 = $signed(T11746) / $signed(22'h100000);
  assign T11746 = $signed(31'h2b451a54) * $signed(16'hffff);
  assign T11747 = $signed(T11748) / $signed(22'h100000);
  assign T11748 = $signed(31'h2f2800ae) * $signed(16'h0);
  assign T11749 = T10817[1'h0:1'h0];
  assign T11750 = T11759 ? twiddle4_2_123_imag : twiddle4_2_122_imag;
  assign twiddle4_2_122_imag = T11753 + T11751;
  assign T11751 = $signed(T11752) / $signed(22'h100000);
  assign T11752 = $signed(31'h2b8ef77c) * $signed(16'hffff);
  assign T11753 = $signed(T11754) / $signed(22'h100000);
  assign T11754 = $signed(31'h2ee3cebe) * $signed(16'h0);
  assign twiddle4_2_123_imag = T11757 + T11755;
  assign T11755 = $signed(T11756) / $signed(22'h100000);
  assign T11756 = $signed(31'h2bd8692b) * $signed(16'hffff);
  assign T11757 = $signed(T11758) / $signed(22'h100000);
  assign T11758 = $signed(31'h2e9f291b) * $signed(16'h0);
  assign T11759 = T10817[1'h0:1'h0];
  assign T11760 = T10817[1'h1:1'h1];
  assign T11761 = T11782 ? T11772 : T11762;
  assign T11762 = T11771 ? twiddle4_2_125_imag : twiddle4_2_124_imag;
  assign twiddle4_2_124_imag = T11765 + T11763;
  assign T11763 = $signed(T11764) / $signed(22'h100000);
  assign T11764 = $signed(31'h2c216eaa) * $signed(16'hffff);
  assign T11765 = $signed(T11766) / $signed(22'h100000);
  assign T11766 = $signed(31'h2e5a106f) * $signed(16'h0);
  assign twiddle4_2_125_imag = T11769 + T11767;
  assign T11767 = $signed(T11768) / $signed(22'h100000);
  assign T11768 = $signed(31'h2c6a0746) * $signed(16'hffff);
  assign T11769 = $signed(T11770) / $signed(22'h100000);
  assign T11770 = $signed(31'h2e148566) * $signed(16'h0);
  assign T11771 = T10817[1'h0:1'h0];
  assign T11772 = T11781 ? twiddle4_2_127_imag : twiddle4_2_126_imag;
  assign twiddle4_2_126_imag = T11775 + T11773;
  assign T11773 = $signed(T11774) / $signed(22'h100000);
  assign T11774 = $signed(31'h2cb2324b) * $signed(16'hffff);
  assign T11775 = $signed(T11776) / $signed(22'h100000);
  assign T11776 = $signed(31'h2dce88a9) * $signed(16'h0);
  assign twiddle4_2_127_imag = T11779 + T11777;
  assign T11777 = $signed(T11778) / $signed(22'h100000);
  assign T11778 = $signed(31'h2cf9ef09) * $signed(16'hffff);
  assign T11779 = $signed(T11780) / $signed(22'h100000);
  assign T11780 = $signed(31'h2d881ae7) * $signed(16'h0);
  assign T11781 = T10817[1'h0:1'h0];
  assign T11782 = T10817[1'h1:1'h1];
  assign T11783 = T10817[2'h2:2'h2];
  assign T11784 = T10817[2'h3:2'h3];
  assign T11785 = T10817[3'h4:3'h4];
  assign T11786 = T10817[3'h5:3'h5];
  assign T11787 = T11361[6'h2e:6'h2e];
  assign T11788 = T10817[3'h6:3'h6];
  assign T11789 = {T12767, T11790};
  assign T11790 = T12766 ? T12215 : T11791;
  assign T11791 = T12214 ? T11982 : T11792;
  assign T11792 = T11981 ? T11887 : T11793;
  assign T11793 = T11886 ? T11840 : T11794;
  assign T11794 = T11839 ? T11817 : T11795;
  assign T11795 = T11816 ? T11806 : T11796;
  assign T11796 = T11805 ? twiddle4_2_129_imag : twiddle4_2_128_imag;
  assign twiddle4_2_128_imag = T11799 + T11797;
  assign T11797 = $signed(T11798) / $signed(22'h100000);
  assign T11798 = $signed(31'h2d413ccc) * $signed(16'hffff);
  assign T11799 = $signed(T11800) / $signed(22'h100000);
  assign T11800 = $signed(31'h2d413ccc) * $signed(16'h0);
  assign twiddle4_2_129_imag = T11803 + T11801;
  assign T11801 = $signed(T11802) / $signed(22'h100000);
  assign T11802 = $signed(31'h2d881ae7) * $signed(16'hffff);
  assign T11803 = $signed(T11804) / $signed(22'h100000);
  assign T11804 = $signed(31'h2cf9ef09) * $signed(16'h0);
  assign T11805 = T10817[1'h0:1'h0];
  assign T11806 = T11815 ? twiddle4_2_131_imag : twiddle4_2_130_imag;
  assign twiddle4_2_130_imag = T11809 + T11807;
  assign T11807 = $signed(T11808) / $signed(22'h100000);
  assign T11808 = $signed(31'h2dce88a9) * $signed(16'hffff);
  assign T11809 = $signed(T11810) / $signed(22'h100000);
  assign T11810 = $signed(31'h2cb2324b) * $signed(16'h0);
  assign twiddle4_2_131_imag = T11813 + T11811;
  assign T11811 = $signed(T11812) / $signed(22'h100000);
  assign T11812 = $signed(31'h2e148566) * $signed(16'hffff);
  assign T11813 = $signed(T11814) / $signed(22'h100000);
  assign T11814 = $signed(31'h2c6a0746) * $signed(16'h0);
  assign T11815 = T10817[1'h0:1'h0];
  assign T11816 = T10817[1'h1:1'h1];
  assign T11817 = T11838 ? T11828 : T11818;
  assign T11818 = T11827 ? twiddle4_2_133_imag : twiddle4_2_132_imag;
  assign twiddle4_2_132_imag = T11821 + T11819;
  assign T11819 = $signed(T11820) / $signed(22'h100000);
  assign T11820 = $signed(31'h2e5a106f) * $signed(16'hffff);
  assign T11821 = $signed(T11822) / $signed(22'h100000);
  assign T11822 = $signed(31'h2c216eaa) * $signed(16'h0);
  assign twiddle4_2_133_imag = T11825 + T11823;
  assign T11823 = $signed(T11824) / $signed(22'h100000);
  assign T11824 = $signed(31'h2e9f291b) * $signed(16'hffff);
  assign T11825 = $signed(T11826) / $signed(22'h100000);
  assign T11826 = $signed(31'h2bd8692b) * $signed(16'h0);
  assign T11827 = T10817[1'h0:1'h0];
  assign T11828 = T11837 ? twiddle4_2_135_imag : twiddle4_2_134_imag;
  assign twiddle4_2_134_imag = T11831 + T11829;
  assign T11829 = $signed(T11830) / $signed(22'h100000);
  assign T11830 = $signed(31'h2ee3cebe) * $signed(16'hffff);
  assign T11831 = $signed(T11832) / $signed(22'h100000);
  assign T11832 = $signed(31'h2b8ef77c) * $signed(16'h0);
  assign twiddle4_2_135_imag = T11835 + T11833;
  assign T11833 = $signed(T11834) / $signed(22'h100000);
  assign T11834 = $signed(31'h2f2800ae) * $signed(16'hffff);
  assign T11835 = $signed(T11836) / $signed(22'h100000);
  assign T11836 = $signed(31'h2b451a54) * $signed(16'h0);
  assign T11837 = T10817[1'h0:1'h0];
  assign T11838 = T10817[1'h1:1'h1];
  assign T11839 = T10817[2'h2:2'h2];
  assign T11840 = T11885 ? T11863 : T11841;
  assign T11841 = T11862 ? T11852 : T11842;
  assign T11842 = T11851 ? twiddle4_2_137_imag : twiddle4_2_136_imag;
  assign twiddle4_2_136_imag = T11845 + T11843;
  assign T11843 = $signed(T11844) / $signed(22'h100000);
  assign T11844 = $signed(31'h2f6bbe44) * $signed(16'hffff);
  assign T11845 = $signed(T11846) / $signed(22'h100000);
  assign T11846 = $signed(31'h2afad269) * $signed(16'h0);
  assign twiddle4_2_137_imag = T11849 + T11847;
  assign T11847 = $signed(T11848) / $signed(22'h100000);
  assign T11848 = $signed(31'h2faf06d9) * $signed(16'hffff);
  assign T11849 = $signed(T11850) / $signed(22'h100000);
  assign T11850 = $signed(31'h2ab02071) * $signed(16'h0);
  assign T11851 = T10817[1'h0:1'h0];
  assign T11852 = T11861 ? twiddle4_2_139_imag : twiddle4_2_138_imag;
  assign twiddle4_2_138_imag = T11855 + T11853;
  assign T11853 = $signed(T11854) / $signed(22'h100000);
  assign T11854 = $signed(31'h2ff1d9c6) * $signed(16'hffff);
  assign T11855 = $signed(T11856) / $signed(22'h100000);
  assign T11856 = $signed(31'h2a650525) * $signed(16'h0);
  assign twiddle4_2_139_imag = T11859 + T11857;
  assign T11857 = $signed(T11858) / $signed(22'h100000);
  assign T11858 = $signed(31'h30343667) * $signed(16'hffff);
  assign T11859 = $signed(T11860) / $signed(22'h100000);
  assign T11860 = $signed(31'h2a19813e) * $signed(16'h0);
  assign T11861 = T10817[1'h0:1'h0];
  assign T11862 = T10817[1'h1:1'h1];
  assign T11863 = T11884 ? T11874 : T11864;
  assign T11864 = T11873 ? twiddle4_2_141_imag : twiddle4_2_140_imag;
  assign twiddle4_2_140_imag = T11867 + T11865;
  assign T11865 = $signed(T11866) / $signed(22'h100000);
  assign T11866 = $signed(31'h30761c17) * $signed(16'hffff);
  assign T11867 = $signed(T11868) / $signed(22'h100000);
  assign T11868 = $signed(31'h29cd9577) * $signed(16'h0);
  assign twiddle4_2_141_imag = T11871 + T11869;
  assign T11869 = $signed(T11870) / $signed(22'h100000);
  assign T11870 = $signed(31'h30b78a35) * $signed(16'hffff);
  assign T11871 = $signed(T11872) / $signed(22'h100000);
  assign T11872 = $signed(31'h2981428b) * $signed(16'h0);
  assign T11873 = T10817[1'h0:1'h0];
  assign T11874 = T11883 ? twiddle4_2_143_imag : twiddle4_2_142_imag;
  assign twiddle4_2_142_imag = T11877 + T11875;
  assign T11875 = $signed(T11876) / $signed(22'h100000);
  assign T11876 = $signed(31'h30f8801f) * $signed(16'hffff);
  assign T11877 = $signed(T11878) / $signed(22'h100000);
  assign T11878 = $signed(31'h29348937) * $signed(16'h0);
  assign twiddle4_2_143_imag = T11881 + T11879;
  assign T11879 = $signed(T11880) / $signed(22'h100000);
  assign T11880 = $signed(31'h3138fd34) * $signed(16'hffff);
  assign T11881 = $signed(T11882) / $signed(22'h100000);
  assign T11882 = $signed(31'h28e76a37) * $signed(16'h0);
  assign T11883 = T10817[1'h0:1'h0];
  assign T11884 = T10817[1'h1:1'h1];
  assign T11885 = T10817[2'h2:2'h2];
  assign T11886 = T10817[2'h3:2'h3];
  assign T11887 = T11980 ? T11934 : T11888;
  assign T11888 = T11933 ? T11911 : T11889;
  assign T11889 = T11910 ? T11900 : T11890;
  assign T11890 = T11899 ? twiddle4_2_145_imag : twiddle4_2_144_imag;
  assign twiddle4_2_144_imag = T11893 + T11891;
  assign T11891 = $signed(T11892) / $signed(22'h100000);
  assign T11892 = $signed(31'h317900d6) * $signed(16'hffff);
  assign T11893 = $signed(T11894) / $signed(22'h100000);
  assign T11894 = $signed(31'h2899e64a) * $signed(16'h0);
  assign twiddle4_2_145_imag = T11897 + T11895;
  assign T11895 = $signed(T11896) / $signed(22'h100000);
  assign T11896 = $signed(31'h31b88a66) * $signed(16'hffff);
  assign T11897 = $signed(T11898) / $signed(22'h100000);
  assign T11898 = $signed(31'h284bfe2f) * $signed(16'h0);
  assign T11899 = T10817[1'h0:1'h0];
  assign T11900 = T11909 ? twiddle4_2_147_imag : twiddle4_2_146_imag;
  assign twiddle4_2_146_imag = T11903 + T11901;
  assign T11901 = $signed(T11902) / $signed(22'h100000);
  assign T11902 = $signed(31'h31f79947) * $signed(16'hffff);
  assign T11903 = $signed(T11904) / $signed(22'h100000);
  assign T11904 = $signed(31'h27fdb2a6) * $signed(16'h0);
  assign twiddle4_2_147_imag = T11907 + T11905;
  assign T11905 = $signed(T11906) / $signed(22'h100000);
  assign T11906 = $signed(31'h32362cdf) * $signed(16'hffff);
  assign T11907 = $signed(T11908) / $signed(22'h100000);
  assign T11908 = $signed(31'h27af0471) * $signed(16'h0);
  assign T11909 = T10817[1'h0:1'h0];
  assign T11910 = T10817[1'h1:1'h1];
  assign T11911 = T11932 ? T11922 : T11912;
  assign T11912 = T11921 ? twiddle4_2_149_imag : twiddle4_2_148_imag;
  assign twiddle4_2_148_imag = T11915 + T11913;
  assign T11913 = $signed(T11914) / $signed(22'h100000);
  assign T11914 = $signed(31'h32744493) * $signed(16'hffff);
  assign T11915 = $signed(T11916) / $signed(22'h100000);
  assign T11916 = $signed(31'h275ff452) * $signed(16'h0);
  assign twiddle4_2_149_imag = T11919 + T11917;
  assign T11917 = $signed(T11918) / $signed(22'h100000);
  assign T11918 = $signed(31'h32b1dfc9) * $signed(16'hffff);
  assign T11919 = $signed(T11920) / $signed(22'h100000);
  assign T11920 = $signed(31'h2710830b) * $signed(16'h0);
  assign T11921 = T10817[1'h0:1'h0];
  assign T11922 = T11931 ? twiddle4_2_151_imag : twiddle4_2_150_imag;
  assign twiddle4_2_150_imag = T11925 + T11923;
  assign T11923 = $signed(T11924) / $signed(22'h100000);
  assign T11924 = $signed(31'h32eefde9) * $signed(16'hffff);
  assign T11925 = $signed(T11926) / $signed(22'h100000);
  assign T11926 = $signed(31'h26c0b162) * $signed(16'h0);
  assign twiddle4_2_151_imag = T11929 + T11927;
  assign T11927 = $signed(T11928) / $signed(22'h100000);
  assign T11928 = $signed(31'h332b9e5d) * $signed(16'hffff);
  assign T11929 = $signed(T11930) / $signed(22'h100000);
  assign T11930 = $signed(31'h2670801a) * $signed(16'h0);
  assign T11931 = T10817[1'h0:1'h0];
  assign T11932 = T10817[1'h1:1'h1];
  assign T11933 = T10817[2'h2:2'h2];
  assign T11934 = T11979 ? T11957 : T11935;
  assign T11935 = T11956 ? T11946 : T11936;
  assign T11936 = T11945 ? twiddle4_2_153_imag : twiddle4_2_152_imag;
  assign twiddle4_2_152_imag = T11939 + T11937;
  assign T11937 = $signed(T11938) / $signed(22'h100000);
  assign T11938 = $signed(31'h3367c08f) * $signed(16'hffff);
  assign T11939 = $signed(T11940) / $signed(22'h100000);
  assign T11940 = $signed(31'h261feff9) * $signed(16'h0);
  assign twiddle4_2_153_imag = T11943 + T11941;
  assign T11941 = $signed(T11942) / $signed(22'h100000);
  assign T11942 = $signed(31'h33a363eb) * $signed(16'hffff);
  assign T11943 = $signed(T11944) / $signed(22'h100000);
  assign T11944 = $signed(31'h25cf01c7) * $signed(16'h0);
  assign T11945 = T10817[1'h0:1'h0];
  assign T11946 = T11955 ? twiddle4_2_155_imag : twiddle4_2_154_imag;
  assign twiddle4_2_154_imag = T11949 + T11947;
  assign T11947 = $signed(T11948) / $signed(22'h100000);
  assign T11948 = $signed(31'h33de87de) * $signed(16'hffff);
  assign T11949 = $signed(T11950) / $signed(22'h100000);
  assign T11950 = $signed(31'h257db64b) * $signed(16'h0);
  assign twiddle4_2_155_imag = T11953 + T11951;
  assign T11951 = $signed(T11952) / $signed(22'h100000);
  assign T11952 = $signed(31'h34192bd5) * $signed(16'hffff);
  assign T11953 = $signed(T11954) / $signed(22'h100000);
  assign T11954 = $signed(31'h252c0e4e) * $signed(16'h0);
  assign T11955 = T10817[1'h0:1'h0];
  assign T11956 = T10817[1'h1:1'h1];
  assign T11957 = T11978 ? T11968 : T11958;
  assign T11958 = T11967 ? twiddle4_2_157_imag : twiddle4_2_156_imag;
  assign twiddle4_2_156_imag = T11961 + T11959;
  assign T11959 = $signed(T11960) / $signed(22'h100000);
  assign T11960 = $signed(31'h34534f40) * $signed(16'hffff);
  assign T11961 = $signed(T11962) / $signed(22'h100000);
  assign T11962 = $signed(31'h24da0a99) * $signed(16'h0);
  assign twiddle4_2_157_imag = T11965 + T11963;
  assign T11963 = $signed(T11964) / $signed(22'h100000);
  assign T11964 = $signed(31'h348cf190) * $signed(16'hffff);
  assign T11965 = $signed(T11966) / $signed(22'h100000);
  assign T11966 = $signed(31'h2487abf7) * $signed(16'h0);
  assign T11967 = T10817[1'h0:1'h0];
  assign T11968 = T11977 ? twiddle4_2_159_imag : twiddle4_2_158_imag;
  assign twiddle4_2_158_imag = T11971 + T11969;
  assign T11969 = $signed(T11970) / $signed(22'h100000);
  assign T11970 = $signed(31'h34c61236) * $signed(16'hffff);
  assign T11971 = $signed(T11972) / $signed(22'h100000);
  assign T11972 = $signed(31'h2434f332) * $signed(16'h0);
  assign twiddle4_2_159_imag = T11975 + T11973;
  assign T11973 = $signed(T11974) / $signed(22'h100000);
  assign T11974 = $signed(31'h34feb0a5) * $signed(16'hffff);
  assign T11975 = $signed(T11976) / $signed(22'h100000);
  assign T11976 = $signed(31'h23e1e117) * $signed(16'h0);
  assign T11977 = T10817[1'h0:1'h0];
  assign T11978 = T10817[1'h1:1'h1];
  assign T11979 = T10817[2'h2:2'h2];
  assign T11980 = T10817[2'h3:2'h3];
  assign T11981 = T10817[3'h4:3'h4];
  assign T11982 = T12213 ? T12087 : T11983;
  assign T11983 = T12086 ? T12030 : T11984;
  assign T11984 = T12029 ? T12007 : T11985;
  assign T11985 = T12006 ? T11996 : T11986;
  assign T11986 = T11995 ? twiddle4_2_161_imag : twiddle4_2_160_imag;
  assign twiddle4_2_160_imag = T11989 + T11987;
  assign T11987 = $signed(T11988) / $signed(22'h100000);
  assign T11988 = $signed(31'h3536cc52) * $signed(16'hffff);
  assign T11989 = $signed(T11990) / $signed(22'h100000);
  assign T11990 = $signed(31'h238e7673) * $signed(16'h0);
  assign twiddle4_2_161_imag = T11993 + T11991;
  assign T11991 = $signed(T11992) / $signed(22'h100000);
  assign T11992 = $signed(31'h356e64b2) * $signed(16'hffff);
  assign T11993 = $signed(T11994) / $signed(22'h100000);
  assign T11994 = $signed(31'h233ab413) * $signed(16'h0);
  assign T11995 = T10817[1'h0:1'h0];
  assign T11996 = T12005 ? twiddle4_2_163_imag : twiddle4_2_162_imag;
  assign twiddle4_2_162_imag = T11999 + T11997;
  assign T11997 = $signed(T11998) / $signed(22'h100000);
  assign T11998 = $signed(31'h35a5793c) * $signed(16'hffff);
  assign T11999 = $signed(T12000) / $signed(22'h100000);
  assign T12000 = $signed(31'h22e69ac7) * $signed(16'h0);
  assign twiddle4_2_163_imag = T12003 + T12001;
  assign T12001 = $signed(T12002) / $signed(22'h100000);
  assign T12002 = $signed(31'h35dc0968) * $signed(16'hffff);
  assign T12003 = $signed(T12004) / $signed(22'h100000);
  assign T12004 = $signed(31'h22922b5e) * $signed(16'h0);
  assign T12005 = T10817[1'h0:1'h0];
  assign T12006 = T10817[1'h1:1'h1];
  assign T12007 = T12028 ? T12018 : T12008;
  assign T12008 = T12017 ? twiddle4_2_165_imag : twiddle4_2_164_imag;
  assign twiddle4_2_164_imag = T12011 + T12009;
  assign T12009 = $signed(T12010) / $signed(22'h100000);
  assign T12010 = $signed(31'h361214b0) * $signed(16'hffff);
  assign T12011 = $signed(T12012) / $signed(22'h100000);
  assign T12012 = $signed(31'h223d66a8) * $signed(16'h0);
  assign twiddle4_2_165_imag = T12015 + T12013;
  assign T12013 = $signed(T12014) / $signed(22'h100000);
  assign T12014 = $signed(31'h36479a8e) * $signed(16'hffff);
  assign T12015 = $signed(T12016) / $signed(22'h100000);
  assign T12016 = $signed(31'h21e84d76) * $signed(16'h0);
  assign T12017 = T10817[1'h0:1'h0];
  assign T12018 = T12027 ? twiddle4_2_167_imag : twiddle4_2_166_imag;
  assign twiddle4_2_166_imag = T12021 + T12019;
  assign T12019 = $signed(T12020) / $signed(22'h100000);
  assign T12020 = $signed(31'h367c9a7d) * $signed(16'hffff);
  assign T12021 = $signed(T12022) / $signed(22'h100000);
  assign T12022 = $signed(31'h2192e09a) * $signed(16'h0);
  assign twiddle4_2_167_imag = T12025 + T12023;
  assign T12023 = $signed(T12024) / $signed(22'h100000);
  assign T12024 = $signed(31'h36b113fd) * $signed(16'hffff);
  assign T12025 = $signed(T12026) / $signed(22'h100000);
  assign T12026 = $signed(31'h213d20e8) * $signed(16'h0);
  assign T12027 = T10817[1'h0:1'h0];
  assign T12028 = T10817[1'h1:1'h1];
  assign T12029 = T10817[2'h2:2'h2];
  assign T12030 = T12085 ? T12055 : T12031;
  assign T12031 = T12054 ? T12042 : T12032;
  assign T12032 = T12041 ? twiddle4_2_169_imag : twiddle4_2_168_imag;
  assign twiddle4_2_168_imag = T12035 + T12033;
  assign T12033 = $signed(T12034) / $signed(22'h100000);
  assign T12034 = $signed(31'h36e5068a) * $signed(16'hffff);
  assign T12035 = $signed(T12036) / $signed(22'h100000);
  assign T12036 = $signed(31'h20e70f32) * $signed(16'h0);
  assign twiddle4_2_169_imag = T12039 + T12037;
  assign T12037 = $signed(T12038) / $signed(22'h100000);
  assign T12038 = $signed(31'h371871a4) * $signed(16'hffff);
  assign T12039 = $signed(T12040) / $signed(22'h100000);
  assign T12040 = $signed(31'h2090ac4d) * $signed(16'h0);
  assign T12041 = T10817[1'h0:1'h0];
  assign T12042 = T12053 ? twiddle4_2_171_imag : twiddle4_2_170_imag;
  assign twiddle4_2_170_imag = T12045 + T12043;
  assign T12043 = $signed(T12044) / $signed(22'h100000);
  assign T12044 = $signed(31'h374b54ce) * $signed(16'hffff);
  assign T12045 = $signed(T12046) / $signed(22'h100000);
  assign T12046 = $signed(31'h2039f90e) * $signed(16'h0);
  assign twiddle4_2_171_imag = T12049 + T12047;
  assign T12047 = $signed(T12048) / $signed(22'h100000);
  assign T12048 = $signed(31'h377daf89) * $signed(16'hffff);
  assign T12049 = {T12052, T12050};
  assign T12050 = $signed(T12051) / $signed(22'h100000);
  assign T12051 = $signed(30'h1fe2f64b) * $signed(16'h0);
  assign T12052 = T12050[6'h2d:6'h2d];
  assign T12053 = T10817[1'h0:1'h0];
  assign T12054 = T10817[1'h1:1'h1];
  assign T12055 = T12084 ? T12070 : T12056;
  assign T12056 = T12069 ? twiddle4_2_173_imag : twiddle4_2_172_imag;
  assign twiddle4_2_172_imag = T12059 + T12057;
  assign T12057 = $signed(T12058) / $signed(22'h100000);
  assign T12058 = $signed(31'h37af8158) * $signed(16'hffff);
  assign T12059 = {T12062, T12060};
  assign T12060 = $signed(T12061) / $signed(22'h100000);
  assign T12061 = $signed(30'h1f8ba4db) * $signed(16'h0);
  assign T12062 = T12060[6'h2d:6'h2d];
  assign twiddle4_2_173_imag = T12065 + T12063;
  assign T12063 = $signed(T12064) / $signed(22'h100000);
  assign T12064 = $signed(31'h37e0c9c2) * $signed(16'hffff);
  assign T12065 = {T12068, T12066};
  assign T12066 = $signed(T12067) / $signed(22'h100000);
  assign T12067 = $signed(30'h1f340596) * $signed(16'h0);
  assign T12068 = T12066[6'h2d:6'h2d];
  assign T12069 = T10817[1'h0:1'h0];
  assign T12070 = T12083 ? twiddle4_2_175_imag : twiddle4_2_174_imag;
  assign twiddle4_2_174_imag = T12073 + T12071;
  assign T12071 = $signed(T12072) / $signed(22'h100000);
  assign T12072 = $signed(31'h3811884c) * $signed(16'hffff);
  assign T12073 = {T12076, T12074};
  assign T12074 = $signed(T12075) / $signed(22'h100000);
  assign T12075 = $signed(30'h1edc1952) * $signed(16'h0);
  assign T12076 = T12074[6'h2d:6'h2d];
  assign twiddle4_2_175_imag = T12079 + T12077;
  assign T12077 = $signed(T12078) / $signed(22'h100000);
  assign T12078 = $signed(31'h3841bc7f) * $signed(16'hffff);
  assign T12079 = {T12082, T12080};
  assign T12080 = $signed(T12081) / $signed(22'h100000);
  assign T12081 = $signed(30'h1e83e0ea) * $signed(16'h0);
  assign T12082 = T12080[6'h2d:6'h2d];
  assign T12083 = T10817[1'h0:1'h0];
  assign T12084 = T10817[1'h1:1'h1];
  assign T12085 = T10817[2'h2:2'h2];
  assign T12086 = T10817[2'h3:2'h3];
  assign T12087 = T12212 ? T12150 : T12088;
  assign T12088 = T12149 ? T12119 : T12089;
  assign T12089 = T12118 ? T12104 : T12090;
  assign T12090 = T12103 ? twiddle4_2_177_imag : twiddle4_2_176_imag;
  assign twiddle4_2_176_imag = T12093 + T12091;
  assign T12091 = $signed(T12092) / $signed(22'h100000);
  assign T12092 = $signed(31'h387165e3) * $signed(16'hffff);
  assign T12093 = {T12096, T12094};
  assign T12094 = $signed(T12095) / $signed(22'h100000);
  assign T12095 = $signed(30'h1e2b5d38) * $signed(16'h0);
  assign T12096 = T12094[6'h2d:6'h2d];
  assign twiddle4_2_177_imag = T12099 + T12097;
  assign T12097 = $signed(T12098) / $signed(22'h100000);
  assign T12098 = $signed(31'h38a08402) * $signed(16'hffff);
  assign T12099 = {T12102, T12100};
  assign T12100 = $signed(T12101) / $signed(22'h100000);
  assign T12101 = $signed(30'h1dd28f14) * $signed(16'h0);
  assign T12102 = T12100[6'h2d:6'h2d];
  assign T12103 = T10817[1'h0:1'h0];
  assign T12104 = T12117 ? twiddle4_2_179_imag : twiddle4_2_178_imag;
  assign twiddle4_2_178_imag = T12107 + T12105;
  assign T12105 = $signed(T12106) / $signed(22'h100000);
  assign T12106 = $signed(31'h38cf1669) * $signed(16'hffff);
  assign T12107 = {T12110, T12108};
  assign T12108 = $signed(T12109) / $signed(22'h100000);
  assign T12109 = $signed(30'h1d79775b) * $signed(16'h0);
  assign T12110 = T12108[6'h2d:6'h2d];
  assign twiddle4_2_179_imag = T12113 + T12111;
  assign T12111 = $signed(T12112) / $signed(22'h100000);
  assign T12112 = $signed(31'h38fd1ca4) * $signed(16'hffff);
  assign T12113 = {T12116, T12114};
  assign T12114 = $signed(T12115) / $signed(22'h100000);
  assign T12115 = $signed(30'h1d2016e8) * $signed(16'h0);
  assign T12116 = T12114[6'h2d:6'h2d];
  assign T12117 = T10817[1'h0:1'h0];
  assign T12118 = T10817[1'h1:1'h1];
  assign T12119 = T12148 ? T12134 : T12120;
  assign T12120 = T12133 ? twiddle4_2_181_imag : twiddle4_2_180_imag;
  assign twiddle4_2_180_imag = T12123 + T12121;
  assign T12121 = $signed(T12122) / $signed(22'h100000);
  assign T12122 = $signed(31'h392a9642) * $signed(16'hffff);
  assign T12123 = {T12126, T12124};
  assign T12124 = $signed(T12125) / $signed(22'h100000);
  assign T12125 = $signed(30'h1cc66e99) * $signed(16'h0);
  assign T12126 = T12124[6'h2d:6'h2d];
  assign twiddle4_2_181_imag = T12129 + T12127;
  assign T12127 = $signed(T12128) / $signed(22'h100000);
  assign T12128 = $signed(31'h395782d3) * $signed(16'hffff);
  assign T12129 = {T12132, T12130};
  assign T12130 = $signed(T12131) / $signed(22'h100000);
  assign T12131 = $signed(30'h1c6c7f49) * $signed(16'h0);
  assign T12132 = T12130[6'h2d:6'h2d];
  assign T12133 = T10817[1'h0:1'h0];
  assign T12134 = T12147 ? twiddle4_2_183_imag : twiddle4_2_182_imag;
  assign twiddle4_2_182_imag = T12137 + T12135;
  assign T12135 = $signed(T12136) / $signed(22'h100000);
  assign T12136 = $signed(31'h3983e1e7) * $signed(16'hffff);
  assign T12137 = {T12140, T12138};
  assign T12138 = $signed(T12139) / $signed(22'h100000);
  assign T12139 = $signed(30'h1c1249d8) * $signed(16'h0);
  assign T12140 = T12138[6'h2d:6'h2d];
  assign twiddle4_2_183_imag = T12143 + T12141;
  assign T12141 = $signed(T12142) / $signed(22'h100000);
  assign T12142 = $signed(31'h39afb313) * $signed(16'hffff);
  assign T12143 = {T12146, T12144};
  assign T12144 = $signed(T12145) / $signed(22'h100000);
  assign T12145 = $signed(30'h1bb7cf23) * $signed(16'h0);
  assign T12146 = T12144[6'h2d:6'h2d];
  assign T12147 = T10817[1'h0:1'h0];
  assign T12148 = T10817[1'h1:1'h1];
  assign T12149 = T10817[2'h2:2'h2];
  assign T12150 = T12211 ? T12181 : T12151;
  assign T12151 = T12180 ? T12166 : T12152;
  assign T12152 = T12165 ? twiddle4_2_185_imag : twiddle4_2_184_imag;
  assign twiddle4_2_184_imag = T12155 + T12153;
  assign T12153 = $signed(T12154) / $signed(22'h100000);
  assign T12154 = $signed(31'h39daf5e8) * $signed(16'hffff);
  assign T12155 = {T12158, T12156};
  assign T12156 = $signed(T12157) / $signed(22'h100000);
  assign T12157 = $signed(30'h1b5d1009) * $signed(16'h0);
  assign T12158 = T12156[6'h2d:6'h2d];
  assign twiddle4_2_185_imag = T12161 + T12159;
  assign T12159 = $signed(T12160) / $signed(22'h100000);
  assign T12160 = $signed(31'h3a05a9fd) * $signed(16'hffff);
  assign T12161 = {T12164, T12162};
  assign T12162 = $signed(T12163) / $signed(22'h100000);
  assign T12163 = $signed(30'h1b020d6c) * $signed(16'h0);
  assign T12164 = T12162[6'h2d:6'h2d];
  assign T12165 = T10817[1'h0:1'h0];
  assign T12166 = T12179 ? twiddle4_2_187_imag : twiddle4_2_186_imag;
  assign twiddle4_2_186_imag = T12169 + T12167;
  assign T12167 = $signed(T12168) / $signed(22'h100000);
  assign T12168 = $signed(31'h3a2fcee8) * $signed(16'hffff);
  assign T12169 = {T12172, T12170};
  assign T12170 = $signed(T12171) / $signed(22'h100000);
  assign T12171 = $signed(30'h1aa6c82b) * $signed(16'h0);
  assign T12172 = T12170[6'h2d:6'h2d];
  assign twiddle4_2_187_imag = T12175 + T12173;
  assign T12173 = $signed(T12174) / $signed(22'h100000);
  assign T12174 = $signed(31'h3a596441) * $signed(16'hffff);
  assign T12175 = {T12178, T12176};
  assign T12176 = $signed(T12177) / $signed(22'h100000);
  assign T12177 = $signed(30'h1a4b4127) * $signed(16'h0);
  assign T12178 = T12176[6'h2d:6'h2d];
  assign T12179 = T10817[1'h0:1'h0];
  assign T12180 = T10817[1'h1:1'h1];
  assign T12181 = T12210 ? T12196 : T12182;
  assign T12182 = T12195 ? twiddle4_2_189_imag : twiddle4_2_188_imag;
  assign twiddle4_2_188_imag = T12185 + T12183;
  assign T12183 = $signed(T12184) / $signed(22'h100000);
  assign T12184 = $signed(31'h3a8269a2) * $signed(16'hffff);
  assign T12185 = {T12188, T12186};
  assign T12186 = $signed(T12187) / $signed(22'h100000);
  assign T12187 = $signed(30'h19ef7943) * $signed(16'h0);
  assign T12188 = T12186[6'h2d:6'h2d];
  assign twiddle4_2_189_imag = T12191 + T12189;
  assign T12189 = $signed(T12190) / $signed(22'h100000);
  assign T12190 = $signed(31'h3aaadea5) * $signed(16'hffff);
  assign T12191 = {T12194, T12192};
  assign T12192 = $signed(T12193) / $signed(22'h100000);
  assign T12193 = $signed(30'h19937161) * $signed(16'h0);
  assign T12194 = T12192[6'h2d:6'h2d];
  assign T12195 = T10817[1'h0:1'h0];
  assign T12196 = T12209 ? twiddle4_2_191_imag : twiddle4_2_190_imag;
  assign twiddle4_2_190_imag = T12199 + T12197;
  assign T12197 = $signed(T12198) / $signed(22'h100000);
  assign T12198 = $signed(31'h3ad2c2e7) * $signed(16'hffff);
  assign T12199 = {T12202, T12200};
  assign T12200 = $signed(T12201) / $signed(22'h100000);
  assign T12201 = $signed(30'h19372a63) * $signed(16'h0);
  assign T12202 = T12200[6'h2d:6'h2d];
  assign twiddle4_2_191_imag = T12205 + T12203;
  assign T12203 = $signed(T12204) / $signed(22'h100000);
  assign T12204 = $signed(31'h3afa1605) * $signed(16'hffff);
  assign T12205 = {T12208, T12206};
  assign T12206 = $signed(T12207) / $signed(22'h100000);
  assign T12207 = $signed(30'h18daa52e) * $signed(16'h0);
  assign T12208 = T12206[6'h2d:6'h2d];
  assign T12209 = T10817[1'h0:1'h0];
  assign T12210 = T10817[1'h1:1'h1];
  assign T12211 = T10817[2'h2:2'h2];
  assign T12212 = T10817[2'h3:2'h3];
  assign T12213 = T10817[3'h4:3'h4];
  assign T12214 = T10817[3'h5:3'h5];
  assign T12215 = T12765 ? T12479 : T12216;
  assign T12216 = T12478 ? T12343 : T12217;
  assign T12217 = T12342 ? T12280 : T12218;
  assign T12218 = T12279 ? T12249 : T12219;
  assign T12219 = T12248 ? T12234 : T12220;
  assign T12220 = T12233 ? twiddle4_2_193_imag : twiddle4_2_192_imag;
  assign twiddle4_2_192_imag = T12223 + T12221;
  assign T12221 = $signed(T12222) / $signed(22'h100000);
  assign T12222 = $signed(31'h3b20d79e) * $signed(16'hffff);
  assign T12223 = {T12226, T12224};
  assign T12224 = $signed(T12225) / $signed(22'h100000);
  assign T12225 = $signed(30'h187de2a6) * $signed(16'h0);
  assign T12226 = T12224[6'h2d:6'h2d];
  assign twiddle4_2_193_imag = T12229 + T12227;
  assign T12227 = $signed(T12228) / $signed(22'h100000);
  assign T12228 = $signed(31'h3b470752) * $signed(16'hffff);
  assign T12229 = {T12232, T12230};
  assign T12230 = $signed(T12231) / $signed(22'h100000);
  assign T12231 = $signed(30'h1820e3b0) * $signed(16'h0);
  assign T12232 = T12230[6'h2d:6'h2d];
  assign T12233 = T10817[1'h0:1'h0];
  assign T12234 = T12247 ? twiddle4_2_195_imag : twiddle4_2_194_imag;
  assign twiddle4_2_194_imag = T12237 + T12235;
  assign T12235 = $signed(T12236) / $signed(22'h100000);
  assign T12236 = $signed(31'h3b6ca4c4) * $signed(16'hffff);
  assign T12237 = {T12240, T12238};
  assign T12238 = $signed(T12239) / $signed(22'h100000);
  assign T12239 = $signed(30'h17c3a931) * $signed(16'h0);
  assign T12240 = T12238[6'h2d:6'h2d];
  assign twiddle4_2_195_imag = T12243 + T12241;
  assign T12241 = $signed(T12242) / $signed(22'h100000);
  assign T12242 = $signed(31'h3b91af96) * $signed(16'hffff);
  assign T12243 = {T12246, T12244};
  assign T12244 = $signed(T12245) / $signed(22'h100000);
  assign T12245 = $signed(30'h1766340f) * $signed(16'h0);
  assign T12246 = T12244[6'h2d:6'h2d];
  assign T12247 = T10817[1'h0:1'h0];
  assign T12248 = T10817[1'h1:1'h1];
  assign T12249 = T12278 ? T12264 : T12250;
  assign T12250 = T12263 ? twiddle4_2_197_imag : twiddle4_2_196_imag;
  assign twiddle4_2_196_imag = T12253 + T12251;
  assign T12251 = $signed(T12252) / $signed(22'h100000);
  assign T12252 = $signed(31'h3bb6276d) * $signed(16'hffff);
  assign T12253 = {T12256, T12254};
  assign T12254 = $signed(T12255) / $signed(22'h100000);
  assign T12255 = $signed(30'h17088530) * $signed(16'h0);
  assign T12256 = T12254[6'h2d:6'h2d];
  assign twiddle4_2_197_imag = T12259 + T12257;
  assign T12257 = $signed(T12258) / $signed(22'h100000);
  assign T12258 = $signed(31'h3bda0bef) * $signed(16'hffff);
  assign T12259 = {T12262, T12260};
  assign T12260 = $signed(T12261) / $signed(22'h100000);
  assign T12261 = $signed(30'h16aa9d7d) * $signed(16'h0);
  assign T12262 = T12260[6'h2d:6'h2d];
  assign T12263 = T10817[1'h0:1'h0];
  assign T12264 = T12277 ? twiddle4_2_199_imag : twiddle4_2_198_imag;
  assign twiddle4_2_198_imag = T12267 + T12265;
  assign T12265 = $signed(T12266) / $signed(22'h100000);
  assign T12266 = $signed(31'h3bfd5cc4) * $signed(16'hffff);
  assign T12267 = {T12270, T12268};
  assign T12268 = $signed(T12269) / $signed(22'h100000);
  assign T12269 = $signed(30'h164c7ddd) * $signed(16'h0);
  assign T12270 = T12268[6'h2d:6'h2d];
  assign twiddle4_2_199_imag = T12273 + T12271;
  assign T12271 = $signed(T12272) / $signed(22'h100000);
  assign T12272 = $signed(31'h3c201994) * $signed(16'hffff);
  assign T12273 = {T12276, T12274};
  assign T12274 = $signed(T12275) / $signed(22'h100000);
  assign T12275 = $signed(30'h15ee2737) * $signed(16'h0);
  assign T12276 = T12274[6'h2d:6'h2d];
  assign T12277 = T10817[1'h0:1'h0];
  assign T12278 = T10817[1'h1:1'h1];
  assign T12279 = T10817[2'h2:2'h2];
  assign T12280 = T12341 ? T12311 : T12281;
  assign T12281 = T12310 ? T12296 : T12282;
  assign T12282 = T12295 ? twiddle4_2_201_imag : twiddle4_2_200_imag;
  assign twiddle4_2_200_imag = T12285 + T12283;
  assign T12283 = $signed(T12284) / $signed(22'h100000);
  assign T12284 = $signed(31'h3c424209) * $signed(16'hffff);
  assign T12285 = {T12288, T12286};
  assign T12286 = $signed(T12287) / $signed(22'h100000);
  assign T12287 = $signed(30'h158f9a75) * $signed(16'h0);
  assign T12288 = T12286[6'h2d:6'h2d];
  assign twiddle4_2_201_imag = T12291 + T12289;
  assign T12289 = $signed(T12290) / $signed(22'h100000);
  assign T12290 = $signed(31'h3c63d5d0) * $signed(16'hffff);
  assign T12291 = {T12294, T12292};
  assign T12292 = $signed(T12293) / $signed(22'h100000);
  assign T12293 = $signed(30'h1530d880) * $signed(16'h0);
  assign T12294 = T12292[6'h2d:6'h2d];
  assign T12295 = T10817[1'h0:1'h0];
  assign T12296 = T12309 ? twiddle4_2_203_imag : twiddle4_2_202_imag;
  assign twiddle4_2_202_imag = T12299 + T12297;
  assign T12297 = $signed(T12298) / $signed(22'h100000);
  assign T12298 = $signed(31'h3c84d496) * $signed(16'hffff);
  assign T12299 = {T12302, T12300};
  assign T12300 = $signed(T12301) / $signed(22'h100000);
  assign T12301 = $signed(30'h14d1e242) * $signed(16'h0);
  assign T12302 = T12300[6'h2d:6'h2d];
  assign twiddle4_2_203_imag = T12305 + T12303;
  assign T12303 = $signed(T12304) / $signed(22'h100000);
  assign T12304 = $signed(31'h3ca53e08) * $signed(16'hffff);
  assign T12305 = {T12308, T12306};
  assign T12306 = $signed(T12307) / $signed(22'h100000);
  assign T12307 = $signed(30'h1472b8a5) * $signed(16'h0);
  assign T12308 = T12306[6'h2d:6'h2d];
  assign T12309 = T10817[1'h0:1'h0];
  assign T12310 = T10817[1'h1:1'h1];
  assign T12311 = T12340 ? T12326 : T12312;
  assign T12312 = T12325 ? twiddle4_2_205_imag : twiddle4_2_204_imag;
  assign twiddle4_2_204_imag = T12315 + T12313;
  assign T12313 = $signed(T12314) / $signed(22'h100000);
  assign T12314 = $signed(31'h3cc511d8) * $signed(16'hffff);
  assign T12315 = {T12318, T12316};
  assign T12316 = $signed(T12317) / $signed(22'h100000);
  assign T12317 = $signed(30'h14135c94) * $signed(16'h0);
  assign T12318 = T12316[6'h2d:6'h2d];
  assign twiddle4_2_205_imag = T12321 + T12319;
  assign T12319 = $signed(T12320) / $signed(22'h100000);
  assign T12320 = $signed(31'h3ce44fb6) * $signed(16'hffff);
  assign T12321 = {T12324, T12322};
  assign T12322 = $signed(T12323) / $signed(22'h100000);
  assign T12323 = $signed(30'h13b3cefa) * $signed(16'h0);
  assign T12324 = T12322[6'h2d:6'h2d];
  assign T12325 = T10817[1'h0:1'h0];
  assign T12326 = T12339 ? twiddle4_2_207_imag : twiddle4_2_206_imag;
  assign twiddle4_2_206_imag = T12329 + T12327;
  assign T12327 = $signed(T12328) / $signed(22'h100000);
  assign T12328 = $signed(31'h3d02f756) * $signed(16'hffff);
  assign T12329 = {T12332, T12330};
  assign T12330 = $signed(T12331) / $signed(22'h100000);
  assign T12331 = $signed(30'h135410c2) * $signed(16'h0);
  assign T12332 = T12330[6'h2d:6'h2d];
  assign twiddle4_2_207_imag = T12335 + T12333;
  assign T12333 = $signed(T12334) / $signed(22'h100000);
  assign T12334 = $signed(31'h3d21086c) * $signed(16'hffff);
  assign T12335 = {T12338, T12336};
  assign T12336 = $signed(T12337) / $signed(22'h100000);
  assign T12337 = $signed(30'h12f422da) * $signed(16'h0);
  assign T12338 = T12336[6'h2d:6'h2d];
  assign T12339 = T10817[1'h0:1'h0];
  assign T12340 = T10817[1'h1:1'h1];
  assign T12341 = T10817[2'h2:2'h2];
  assign T12342 = T10817[2'h3:2'h3];
  assign T12343 = T12477 ? T12407 : T12344;
  assign T12344 = T12406 ? T12375 : T12345;
  assign T12345 = T12374 ? T12360 : T12346;
  assign T12346 = T12359 ? twiddle4_2_209_imag : twiddle4_2_208_imag;
  assign twiddle4_2_208_imag = T12349 + T12347;
  assign T12347 = $signed(T12348) / $signed(22'h100000);
  assign T12348 = $signed(31'h3d3e82ad) * $signed(16'hffff);
  assign T12349 = {T12352, T12350};
  assign T12350 = $signed(T12351) / $signed(22'h100000);
  assign T12351 = $signed(30'h1294062e) * $signed(16'h0);
  assign T12352 = T12350[6'h2d:6'h2d];
  assign twiddle4_2_209_imag = T12355 + T12353;
  assign T12353 = $signed(T12354) / $signed(22'h100000);
  assign T12354 = $signed(31'h3d5b65d1) * $signed(16'hffff);
  assign T12355 = {T12358, T12356};
  assign T12356 = $signed(T12357) / $signed(22'h100000);
  assign T12357 = $signed(30'h1233bbab) * $signed(16'h0);
  assign T12358 = T12356[6'h2d:6'h2d];
  assign T12359 = T10817[1'h0:1'h0];
  assign T12360 = T12373 ? twiddle4_2_211_imag : twiddle4_2_210_imag;
  assign twiddle4_2_210_imag = T12363 + T12361;
  assign T12361 = $signed(T12362) / $signed(22'h100000);
  assign T12362 = $signed(31'h3d77b191) * $signed(16'hffff);
  assign T12363 = {T12366, T12364};
  assign T12364 = $signed(T12365) / $signed(22'h100000);
  assign T12365 = $signed(30'h11d3443f) * $signed(16'h0);
  assign T12366 = T12364[6'h2d:6'h2d];
  assign twiddle4_2_211_imag = T12369 + T12367;
  assign T12367 = $signed(T12368) / $signed(22'h100000);
  assign T12368 = $signed(31'h3d9365a7) * $signed(16'hffff);
  assign T12369 = {T12372, T12370};
  assign T12370 = $signed(T12371) / $signed(22'h100000);
  assign T12371 = $signed(30'h1172a0d7) * $signed(16'h0);
  assign T12372 = T12370[6'h2d:6'h2d];
  assign T12373 = T10817[1'h0:1'h0];
  assign T12374 = T10817[1'h1:1'h1];
  assign T12375 = T12405 ? T12390 : T12376;
  assign T12376 = T12389 ? twiddle4_2_213_imag : twiddle4_2_212_imag;
  assign twiddle4_2_212_imag = T12379 + T12377;
  assign T12377 = $signed(T12378) / $signed(22'h100000);
  assign T12378 = $signed(31'h3dae81ce) * $signed(16'hffff);
  assign T12379 = {T12382, T12380};
  assign T12380 = $signed(T12381) / $signed(22'h100000);
  assign T12381 = $signed(30'h1111d262) * $signed(16'h0);
  assign T12382 = T12380[6'h2d:6'h2d];
  assign twiddle4_2_213_imag = T12385 + T12383;
  assign T12383 = $signed(T12384) / $signed(22'h100000);
  assign T12384 = $signed(31'h3dc905c4) * $signed(16'hffff);
  assign T12385 = {T12388, T12386};
  assign T12386 = $signed(T12387) / $signed(22'h100000);
  assign T12387 = $signed(30'h10b0d9cf) * $signed(16'h0);
  assign T12388 = T12386[6'h2d:6'h2d];
  assign T12389 = T10817[1'h0:1'h0];
  assign T12390 = T12404 ? twiddle4_2_215_imag : twiddle4_2_214_imag;
  assign twiddle4_2_214_imag = T12393 + T12391;
  assign T12391 = $signed(T12392) / $signed(22'h100000);
  assign T12392 = $signed(31'h3de2f147) * $signed(16'hffff);
  assign T12393 = {T12396, T12394};
  assign T12394 = $signed(T12395) / $signed(22'h100000);
  assign T12395 = $signed(30'h104fb80e) * $signed(16'h0);
  assign T12396 = T12394[6'h2d:6'h2d];
  assign twiddle4_2_215_imag = T12399 + T12397;
  assign T12397 = $signed(T12398) / $signed(22'h100000);
  assign T12398 = $signed(31'h3dfc4418) * $signed(16'hffff);
  assign T12399 = {T12402, T12400};
  assign T12400 = $signed(T12401) / $signed(22'h100000);
  assign T12401 = $signed(29'hfee6e0d) * $signed(16'h0);
  assign T12402 = T12403 ? 2'h3 : 2'h0;
  assign T12403 = T12400[6'h2c:6'h2c];
  assign T12404 = T10817[1'h0:1'h0];
  assign T12405 = T10817[1'h1:1'h1];
  assign T12406 = T10817[2'h2:2'h2];
  assign T12407 = T12476 ? T12442 : T12408;
  assign T12408 = T12441 ? T12425 : T12409;
  assign T12409 = T12424 ? twiddle4_2_217_imag : twiddle4_2_216_imag;
  assign twiddle4_2_216_imag = T12412 + T12410;
  assign T12410 = $signed(T12411) / $signed(22'h100000);
  assign T12411 = $signed(31'h3e14fdf7) * $signed(16'hffff);
  assign T12412 = {T12415, T12413};
  assign T12413 = $signed(T12414) / $signed(22'h100000);
  assign T12414 = $signed(29'hf8cfcbd) * $signed(16'h0);
  assign T12415 = T12416 ? 2'h3 : 2'h0;
  assign T12416 = T12413[6'h2c:6'h2c];
  assign twiddle4_2_217_imag = T12419 + T12417;
  assign T12417 = $signed(T12418) / $signed(22'h100000);
  assign T12418 = $signed(31'h3e2d1ea7) * $signed(16'hffff);
  assign T12419 = {T12422, T12420};
  assign T12420 = $signed(T12421) / $signed(22'h100000);
  assign T12421 = $signed(29'hf2b650f) * $signed(16'h0);
  assign T12422 = T12423 ? 2'h3 : 2'h0;
  assign T12423 = T12420[6'h2c:6'h2c];
  assign T12424 = T10817[1'h0:1'h0];
  assign T12425 = T12440 ? twiddle4_2_219_imag : twiddle4_2_218_imag;
  assign twiddle4_2_218_imag = T12428 + T12426;
  assign T12426 = $signed(T12427) / $signed(22'h100000);
  assign T12427 = $signed(31'h3e44a5ee) * $signed(16'hffff);
  assign T12428 = {T12431, T12429};
  assign T12429 = $signed(T12430) / $signed(22'h100000);
  assign T12430 = $signed(29'hec9a7f2) * $signed(16'h0);
  assign T12431 = T12432 ? 2'h3 : 2'h0;
  assign T12432 = T12429[6'h2c:6'h2c];
  assign twiddle4_2_219_imag = T12435 + T12433;
  assign T12433 = $signed(T12434) / $signed(22'h100000);
  assign T12434 = $signed(31'h3e5b9392) * $signed(16'hffff);
  assign T12435 = {T12438, T12436};
  assign T12436 = $signed(T12437) / $signed(22'h100000);
  assign T12437 = $signed(29'he67c659) * $signed(16'h0);
  assign T12438 = T12439 ? 2'h3 : 2'h0;
  assign T12439 = T12436[6'h2c:6'h2c];
  assign T12440 = T10817[1'h0:1'h0];
  assign T12441 = T10817[1'h1:1'h1];
  assign T12442 = T12475 ? T12459 : T12443;
  assign T12443 = T12458 ? twiddle4_2_221_imag : twiddle4_2_220_imag;
  assign twiddle4_2_220_imag = T12446 + T12444;
  assign T12444 = $signed(T12445) / $signed(22'h100000);
  assign T12445 = $signed(31'h3e71e758) * $signed(16'hffff);
  assign T12446 = {T12449, T12447};
  assign T12447 = $signed(T12448) / $signed(22'h100000);
  assign T12448 = $signed(29'he05c135) * $signed(16'h0);
  assign T12449 = T12450 ? 2'h3 : 2'h0;
  assign T12450 = T12447[6'h2c:6'h2c];
  assign twiddle4_2_221_imag = T12453 + T12451;
  assign T12451 = $signed(T12452) / $signed(22'h100000);
  assign T12452 = $signed(31'h3e87a10b) * $signed(16'hffff);
  assign T12453 = {T12456, T12454};
  assign T12454 = $signed(T12455) / $signed(22'h100000);
  assign T12455 = $signed(29'hda39977) * $signed(16'h0);
  assign T12456 = T12457 ? 2'h3 : 2'h0;
  assign T12457 = T12454[6'h2c:6'h2c];
  assign T12458 = T10817[1'h0:1'h0];
  assign T12459 = T12474 ? twiddle4_2_223_imag : twiddle4_2_222_imag;
  assign twiddle4_2_222_imag = T12462 + T12460;
  assign T12460 = $signed(T12461) / $signed(22'h100000);
  assign T12461 = $signed(31'h3e9cc076) * $signed(16'hffff);
  assign T12462 = {T12465, T12463};
  assign T12463 = $signed(T12464) / $signed(22'h100000);
  assign T12464 = $signed(29'hd415012) * $signed(16'h0);
  assign T12465 = T12466 ? 2'h3 : 2'h0;
  assign T12466 = T12463[6'h2c:6'h2c];
  assign twiddle4_2_223_imag = T12469 + T12467;
  assign T12467 = $signed(T12468) / $signed(22'h100000);
  assign T12468 = $signed(31'h3eb14562) * $signed(16'hffff);
  assign T12469 = {T12472, T12470};
  assign T12470 = $signed(T12471) / $signed(22'h100000);
  assign T12471 = $signed(29'hcdee5f9) * $signed(16'h0);
  assign T12472 = T12473 ? 2'h3 : 2'h0;
  assign T12473 = T12470[6'h2c:6'h2c];
  assign T12474 = T10817[1'h0:1'h0];
  assign T12475 = T10817[1'h1:1'h1];
  assign T12476 = T10817[2'h2:2'h2];
  assign T12477 = T10817[2'h3:2'h3];
  assign T12478 = T10817[3'h4:3'h4];
  assign T12479 = T12764 ? T12622 : T12480;
  assign T12480 = T12621 ? T12551 : T12481;
  assign T12481 = T12550 ? T12516 : T12482;
  assign T12482 = T12515 ? T12499 : T12483;
  assign T12483 = T12498 ? twiddle4_2_225_imag : twiddle4_2_224_imag;
  assign twiddle4_2_224_imag = T12486 + T12484;
  assign T12484 = $signed(T12485) / $signed(22'h100000);
  assign T12485 = $signed(31'h3ec52f9f) * $signed(16'hffff);
  assign T12486 = {T12489, T12487};
  assign T12487 = $signed(T12488) / $signed(22'h100000);
  assign T12488 = $signed(29'hc7c5c1e) * $signed(16'h0);
  assign T12489 = T12490 ? 2'h3 : 2'h0;
  assign T12490 = T12487[6'h2c:6'h2c];
  assign twiddle4_2_225_imag = T12493 + T12491;
  assign T12491 = $signed(T12492) / $signed(22'h100000);
  assign T12492 = $signed(31'h3ed87efb) * $signed(16'hffff);
  assign T12493 = {T12496, T12494};
  assign T12494 = $signed(T12495) / $signed(22'h100000);
  assign T12495 = $signed(29'hc19b374) * $signed(16'h0);
  assign T12496 = T12497 ? 2'h3 : 2'h0;
  assign T12497 = T12494[6'h2c:6'h2c];
  assign T12498 = T10817[1'h0:1'h0];
  assign T12499 = T12514 ? twiddle4_2_227_imag : twiddle4_2_226_imag;
  assign twiddle4_2_226_imag = T12502 + T12500;
  assign T12500 = $signed(T12501) / $signed(22'h100000);
  assign T12501 = $signed(31'h3eeb3347) * $signed(16'hffff);
  assign T12502 = {T12505, T12503};
  assign T12503 = $signed(T12504) / $signed(22'h100000);
  assign T12504 = $signed(29'hbb6ecef) * $signed(16'h0);
  assign T12505 = T12506 ? 2'h3 : 2'h0;
  assign T12506 = T12503[6'h2c:6'h2c];
  assign twiddle4_2_227_imag = T12509 + T12507;
  assign T12507 = $signed(T12508) / $signed(22'h100000);
  assign T12508 = $signed(31'h3efd4c53) * $signed(16'hffff);
  assign T12509 = {T12512, T12510};
  assign T12510 = $signed(T12511) / $signed(22'h100000);
  assign T12511 = $signed(29'hb540982) * $signed(16'h0);
  assign T12512 = T12513 ? 2'h3 : 2'h0;
  assign T12513 = T12510[6'h2c:6'h2c];
  assign T12514 = T10817[1'h0:1'h0];
  assign T12515 = T10817[1'h1:1'h1];
  assign T12516 = T12549 ? T12533 : T12517;
  assign T12517 = T12532 ? twiddle4_2_229_imag : twiddle4_2_228_imag;
  assign twiddle4_2_228_imag = T12520 + T12518;
  assign T12518 = $signed(T12519) / $signed(22'h100000);
  assign T12519 = $signed(31'h3f0ec9f4) * $signed(16'hffff);
  assign T12520 = {T12523, T12521};
  assign T12521 = $signed(T12522) / $signed(22'h100000);
  assign T12522 = $signed(29'haf10a22) * $signed(16'h0);
  assign T12523 = T12524 ? 2'h3 : 2'h0;
  assign T12524 = T12521[6'h2c:6'h2c];
  assign twiddle4_2_229_imag = T12527 + T12525;
  assign T12525 = $signed(T12526) / $signed(22'h100000);
  assign T12526 = $signed(31'h3f1fabff) * $signed(16'hffff);
  assign T12527 = {T12530, T12528};
  assign T12528 = $signed(T12529) / $signed(22'h100000);
  assign T12529 = $signed(29'ha8defc2) * $signed(16'h0);
  assign T12530 = T12531 ? 2'h3 : 2'h0;
  assign T12531 = T12528[6'h2c:6'h2c];
  assign T12532 = T10817[1'h0:1'h0];
  assign T12533 = T12548 ? twiddle4_2_231_imag : twiddle4_2_230_imag;
  assign twiddle4_2_230_imag = T12536 + T12534;
  assign T12534 = $signed(T12535) / $signed(22'h100000);
  assign T12535 = $signed(31'h3f2ff249) * $signed(16'hffff);
  assign T12536 = {T12539, T12537};
  assign T12537 = $signed(T12538) / $signed(22'h100000);
  assign T12538 = $signed(29'ha2abb58) * $signed(16'h0);
  assign T12539 = T12540 ? 2'h3 : 2'h0;
  assign T12540 = T12537[6'h2c:6'h2c];
  assign twiddle4_2_231_imag = T12543 + T12541;
  assign T12541 = $signed(T12542) / $signed(22'h100000);
  assign T12542 = $signed(31'h3f3f9cab) * $signed(16'hffff);
  assign T12543 = {T12546, T12544};
  assign T12544 = $signed(T12545) / $signed(22'h100000);
  assign T12545 = $signed(29'h9c76dd8) * $signed(16'h0);
  assign T12546 = T12547 ? 2'h3 : 2'h0;
  assign T12547 = T12544[6'h2c:6'h2c];
  assign T12548 = T10817[1'h0:1'h0];
  assign T12549 = T10817[1'h1:1'h1];
  assign T12550 = T10817[2'h2:2'h2];
  assign T12551 = T12620 ? T12586 : T12552;
  assign T12552 = T12585 ? T12569 : T12553;
  assign T12553 = T12568 ? twiddle4_2_233_imag : twiddle4_2_232_imag;
  assign twiddle4_2_232_imag = T12556 + T12554;
  assign T12554 = $signed(T12555) / $signed(22'h100000);
  assign T12555 = $signed(31'h3f4eaafe) * $signed(16'hffff);
  assign T12556 = {T12559, T12557};
  assign T12557 = $signed(T12558) / $signed(22'h100000);
  assign T12558 = $signed(29'h9640837) * $signed(16'h0);
  assign T12559 = T12560 ? 2'h3 : 2'h0;
  assign T12560 = T12557[6'h2c:6'h2c];
  assign twiddle4_2_233_imag = T12563 + T12561;
  assign T12561 = $signed(T12562) / $signed(22'h100000);
  assign T12562 = $signed(31'h3f5d1d1c) * $signed(16'hffff);
  assign T12563 = {T12566, T12564};
  assign T12564 = $signed(T12565) / $signed(22'h100000);
  assign T12565 = $signed(29'h9008b6a) * $signed(16'h0);
  assign T12566 = T12567 ? 2'h3 : 2'h0;
  assign T12567 = T12564[6'h2c:6'h2c];
  assign T12568 = T10817[1'h0:1'h0];
  assign T12569 = T12584 ? twiddle4_2_235_imag : twiddle4_2_234_imag;
  assign twiddle4_2_234_imag = T12572 + T12570;
  assign T12570 = $signed(T12571) / $signed(22'h100000);
  assign T12571 = $signed(31'h3f6af2e3) * $signed(16'hffff);
  assign T12572 = {T12575, T12573};
  assign T12573 = $signed(T12574) / $signed(22'h100000);
  assign T12574 = $signed(29'h89cf867) * $signed(16'h0);
  assign T12575 = T12576 ? 2'h3 : 2'h0;
  assign T12576 = T12573[6'h2c:6'h2c];
  assign twiddle4_2_235_imag = T12579 + T12577;
  assign T12577 = $signed(T12578) / $signed(22'h100000);
  assign T12578 = $signed(31'h3f782c2f) * $signed(16'hffff);
  assign T12579 = {T12582, T12580};
  assign T12580 = $signed(T12581) / $signed(22'h100000);
  assign T12581 = $signed(29'h8395023) * $signed(16'h0);
  assign T12582 = T12583 ? 2'h3 : 2'h0;
  assign T12583 = T12580[6'h2c:6'h2c];
  assign T12584 = T10817[1'h0:1'h0];
  assign T12585 = T10817[1'h1:1'h1];
  assign T12586 = T12619 ? T12603 : T12587;
  assign T12587 = T12602 ? twiddle4_2_237_imag : twiddle4_2_236_imag;
  assign twiddle4_2_236_imag = T12590 + T12588;
  assign T12588 = $signed(T12589) / $signed(22'h100000);
  assign T12589 = $signed(31'h3f84c8e1) * $signed(16'hffff);
  assign T12590 = {T12593, T12591};
  assign T12591 = $signed(T12592) / $signed(22'h100000);
  assign T12592 = $signed(28'h7d59395) * $signed(16'h0);
  assign T12593 = T12594 ? 3'h7 : 3'h0;
  assign T12594 = T12591[6'h2b:6'h2b];
  assign twiddle4_2_237_imag = T12597 + T12595;
  assign T12595 = $signed(T12596) / $signed(22'h100000);
  assign T12596 = $signed(31'h3f90c8d9) * $signed(16'hffff);
  assign T12597 = {T12600, T12598};
  assign T12598 = $signed(T12599) / $signed(22'h100000);
  assign T12599 = $signed(28'h771c3b2) * $signed(16'h0);
  assign T12600 = T12601 ? 3'h7 : 3'h0;
  assign T12601 = T12598[6'h2b:6'h2b];
  assign T12602 = T10817[1'h0:1'h0];
  assign T12603 = T12618 ? twiddle4_2_239_imag : twiddle4_2_238_imag;
  assign twiddle4_2_238_imag = T12606 + T12604;
  assign T12604 = $signed(T12605) / $signed(22'h100000);
  assign T12605 = $signed(31'h3f9c2bfa) * $signed(16'hffff);
  assign T12606 = {T12609, T12607};
  assign T12607 = $signed(T12608) / $signed(22'h100000);
  assign T12608 = $signed(28'h70de171) * $signed(16'h0);
  assign T12609 = T12610 ? 3'h7 : 3'h0;
  assign T12610 = T12607[6'h2b:6'h2b];
  assign twiddle4_2_239_imag = T12613 + T12611;
  assign T12611 = $signed(T12612) / $signed(22'h100000);
  assign T12612 = $signed(31'h3fa6f228) * $signed(16'hffff);
  assign T12613 = {T12616, T12614};
  assign T12614 = $signed(T12615) / $signed(22'h100000);
  assign T12615 = $signed(28'h6a9edc9) * $signed(16'h0);
  assign T12616 = T12617 ? 3'h7 : 3'h0;
  assign T12617 = T12614[6'h2b:6'h2b];
  assign T12618 = T10817[1'h0:1'h0];
  assign T12619 = T10817[1'h1:1'h1];
  assign T12620 = T10817[2'h2:2'h2];
  assign T12621 = T10817[2'h3:2'h3];
  assign T12622 = T12763 ? T12693 : T12623;
  assign T12623 = T12692 ? T12658 : T12624;
  assign T12624 = T12657 ? T12641 : T12625;
  assign T12625 = T12640 ? twiddle4_2_241_imag : twiddle4_2_240_imag;
  assign twiddle4_2_240_imag = T12628 + T12626;
  assign T12626 = $signed(T12627) / $signed(22'h100000);
  assign T12627 = $signed(31'h3fb11b47) * $signed(16'hffff);
  assign T12628 = {T12631, T12629};
  assign T12629 = $signed(T12630) / $signed(22'h100000);
  assign T12630 = $signed(28'h645e9af) * $signed(16'h0);
  assign T12631 = T12632 ? 3'h7 : 3'h0;
  assign T12632 = T12629[6'h2b:6'h2b];
  assign twiddle4_2_241_imag = T12635 + T12633;
  assign T12633 = $signed(T12634) / $signed(22'h100000);
  assign T12634 = $signed(31'h3fbaa73f) * $signed(16'hffff);
  assign T12635 = {T12638, T12636};
  assign T12636 = $signed(T12637) / $signed(22'h100000);
  assign T12637 = $signed(28'h5e1d61a) * $signed(16'h0);
  assign T12638 = T12639 ? 3'h7 : 3'h0;
  assign T12639 = T12636[6'h2b:6'h2b];
  assign T12640 = T10817[1'h0:1'h0];
  assign T12641 = T12656 ? twiddle4_2_243_imag : twiddle4_2_242_imag;
  assign twiddle4_2_242_imag = T12644 + T12642;
  assign T12642 = $signed(T12643) / $signed(22'h100000);
  assign T12643 = $signed(31'h3fc395f9) * $signed(16'hffff);
  assign T12644 = {T12647, T12645};
  assign T12645 = $signed(T12646) / $signed(22'h100000);
  assign T12646 = $signed(28'h57db402) * $signed(16'h0);
  assign T12647 = T12648 ? 3'h7 : 3'h0;
  assign T12648 = T12645[6'h2b:6'h2b];
  assign twiddle4_2_243_imag = T12651 + T12649;
  assign T12649 = $signed(T12650) / $signed(22'h100000);
  assign T12650 = $signed(31'h3fcbe75e) * $signed(16'hffff);
  assign T12651 = {T12654, T12652};
  assign T12652 = $signed(T12653) / $signed(22'h100000);
  assign T12653 = $signed(28'h519845e) * $signed(16'h0);
  assign T12654 = T12655 ? 3'h7 : 3'h0;
  assign T12655 = T12652[6'h2b:6'h2b];
  assign T12656 = T10817[1'h0:1'h0];
  assign T12657 = T10817[1'h1:1'h1];
  assign T12658 = T12691 ? T12675 : T12659;
  assign T12659 = T12674 ? twiddle4_2_245_imag : twiddle4_2_244_imag;
  assign twiddle4_2_244_imag = T12662 + T12660;
  assign T12660 = $signed(T12661) / $signed(22'h100000);
  assign T12661 = $signed(31'h3fd39b5a) * $signed(16'hffff);
  assign T12662 = {T12665, T12663};
  assign T12663 = $signed(T12664) / $signed(22'h100000);
  assign T12664 = $signed(28'h4b54824) * $signed(16'h0);
  assign T12665 = T12666 ? 3'h7 : 3'h0;
  assign T12666 = T12663[6'h2b:6'h2b];
  assign twiddle4_2_245_imag = T12669 + T12667;
  assign T12667 = $signed(T12668) / $signed(22'h100000);
  assign T12668 = $signed(31'h3fdab1d9) * $signed(16'hffff);
  assign T12669 = {T12672, T12670};
  assign T12670 = $signed(T12671) / $signed(22'h100000);
  assign T12671 = $signed(28'h451004d) * $signed(16'h0);
  assign T12672 = T12673 ? 3'h7 : 3'h0;
  assign T12673 = T12670[6'h2b:6'h2b];
  assign T12674 = T10817[1'h0:1'h0];
  assign T12675 = T12690 ? twiddle4_2_247_imag : twiddle4_2_246_imag;
  assign twiddle4_2_246_imag = T12678 + T12676;
  assign T12676 = $signed(T12677) / $signed(22'h100000);
  assign T12677 = $signed(31'h3fe12acb) * $signed(16'hffff);
  assign T12678 = {T12681, T12679};
  assign T12679 = $signed(T12680) / $signed(22'h100000);
  assign T12680 = $signed(27'h3ecadcf) * $signed(16'h0);
  assign T12681 = T12682 ? 4'hf : 4'h0;
  assign T12682 = T12679[6'h2a:6'h2a];
  assign twiddle4_2_247_imag = T12685 + T12683;
  assign T12683 = $signed(T12684) / $signed(22'h100000);
  assign T12684 = $signed(31'h3fe7061f) * $signed(16'hffff);
  assign T12685 = {T12688, T12686};
  assign T12686 = $signed(T12687) / $signed(22'h100000);
  assign T12687 = $signed(27'h38851a2) * $signed(16'h0);
  assign T12688 = T12689 ? 4'hf : 4'h0;
  assign T12689 = T12686[6'h2a:6'h2a];
  assign T12690 = T10817[1'h0:1'h0];
  assign T12691 = T10817[1'h1:1'h1];
  assign T12692 = T10817[2'h2:2'h2];
  assign T12693 = T12762 ? T12728 : T12694;
  assign T12694 = T12727 ? T12711 : T12695;
  assign T12695 = T12710 ? twiddle4_2_249_imag : twiddle4_2_248_imag;
  assign twiddle4_2_248_imag = T12698 + T12696;
  assign T12696 = $signed(T12697) / $signed(22'h100000);
  assign T12697 = $signed(31'h3fec43c6) * $signed(16'hffff);
  assign T12698 = {T12701, T12699};
  assign T12699 = $signed(T12700) / $signed(22'h100000);
  assign T12700 = $signed(27'h323ecbe) * $signed(16'h0);
  assign T12701 = T12702 ? 4'hf : 4'h0;
  assign T12702 = T12699[6'h2a:6'h2a];
  assign twiddle4_2_249_imag = T12705 + T12703;
  assign T12703 = $signed(T12704) / $signed(22'h100000);
  assign T12704 = $signed(31'h3ff0e3b5) * $signed(16'hffff);
  assign T12705 = {T12708, T12706};
  assign T12706 = $signed(T12707) / $signed(22'h100000);
  assign T12707 = $signed(27'h2bf801a) * $signed(16'h0);
  assign T12708 = T12709 ? 4'hf : 4'h0;
  assign T12709 = T12706[6'h2a:6'h2a];
  assign T12710 = T10817[1'h0:1'h0];
  assign T12711 = T12726 ? twiddle4_2_251_imag : twiddle4_2_250_imag;
  assign twiddle4_2_250_imag = T12714 + T12712;
  assign T12712 = $signed(T12713) / $signed(22'h100000);
  assign T12713 = $signed(31'h3ff4e5df) * $signed(16'hffff);
  assign T12714 = {T12717, T12715};
  assign T12715 = $signed(T12716) / $signed(22'h100000);
  assign T12716 = $signed(27'h25b0cae) * $signed(16'h0);
  assign T12717 = T12718 ? 4'hf : 4'h0;
  assign T12718 = T12715[6'h2a:6'h2a];
  assign twiddle4_2_251_imag = T12721 + T12719;
  assign T12719 = $signed(T12720) / $signed(22'h100000);
  assign T12720 = $signed(31'h3ff84a3b) * $signed(16'hffff);
  assign T12721 = {T12724, T12722};
  assign T12722 = $signed(T12723) / $signed(22'h100000);
  assign T12723 = $signed(26'h1f69373) * $signed(16'h0);
  assign T12724 = T12725 ? 5'h1f : 5'h0;
  assign T12725 = T12722[6'h29:6'h29];
  assign T12726 = T10817[1'h0:1'h0];
  assign T12727 = T10817[1'h1:1'h1];
  assign T12728 = T12761 ? T12745 : T12729;
  assign T12729 = T12744 ? twiddle4_2_253_imag : twiddle4_2_252_imag;
  assign twiddle4_2_252_imag = T12732 + T12730;
  assign T12730 = $signed(T12731) / $signed(22'h100000);
  assign T12731 = $signed(31'h3ffb10c1) * $signed(16'hffff);
  assign T12732 = {T12735, T12733};
  assign T12733 = $signed(T12734) / $signed(22'h100000);
  assign T12734 = $signed(26'h192155f) * $signed(16'h0);
  assign T12735 = T12736 ? 5'h1f : 5'h0;
  assign T12736 = T12733[6'h29:6'h29];
  assign twiddle4_2_253_imag = T12739 + T12737;
  assign T12737 = $signed(T12738) / $signed(22'h100000);
  assign T12738 = $signed(31'h3ffd3968) * $signed(16'hffff);
  assign T12739 = {T12742, T12740};
  assign T12740 = $signed(T12741) / $signed(22'h100000);
  assign T12741 = $signed(26'h12d936b) * $signed(16'h0);
  assign T12742 = T12743 ? 5'h1f : 5'h0;
  assign T12743 = T12740[6'h29:6'h29];
  assign T12744 = T10817[1'h0:1'h0];
  assign T12745 = T12760 ? twiddle4_2_255_imag : twiddle4_2_254_imag;
  assign twiddle4_2_254_imag = T12748 + T12746;
  assign T12746 = $signed(T12747) / $signed(22'h100000);
  assign T12747 = $signed(31'h3ffec42d) * $signed(16'hffff);
  assign T12748 = {T12751, T12749};
  assign T12749 = $signed(T12750) / $signed(22'h100000);
  assign T12750 = $signed(25'hc90e8f) * $signed(16'h0);
  assign T12751 = T12752 ? 6'h3f : 6'h0;
  assign T12752 = T12749[6'h28:6'h28];
  assign twiddle4_2_255_imag = T12755 + T12753;
  assign T12753 = $signed(T12754) / $signed(22'h100000);
  assign T12754 = $signed(31'h3fffb10b) * $signed(16'hffff);
  assign T12755 = {T12758, T12756};
  assign T12756 = $signed(T12757) / $signed(22'h100000);
  assign T12757 = $signed(24'h6487c3) * $signed(16'h0);
  assign T12758 = T12759 ? 7'h7f : 7'h0;
  assign T12759 = T12756[6'h27:6'h27];
  assign T12760 = T10817[1'h0:1'h0];
  assign T12761 = T10817[1'h1:1'h1];
  assign T12762 = T10817[2'h2:2'h2];
  assign T12763 = T10817[2'h3:2'h3];
  assign T12764 = T10817[3'h4:3'h4];
  assign T12765 = T10817[3'h5:3'h5];
  assign T12766 = T10817[3'h6:3'h6];
  assign T12767 = T11790[6'h2e:6'h2e];
  assign T12768 = T10817[3'h7:3'h7];
  assign T12769 = T14743 ? T13764 : T12770;
  assign T12770 = T13763 ? T13335 : T12771;
  assign T12771 = T13334 ? T13068 : T12772;
  assign T12772 = T13067 ? T12923 : T12773;
  assign T12773 = T12922 ? T12850 : T12774;
  assign T12774 = T12849 ? T12813 : T12775;
  assign T12775 = T12812 ? T12794 : T12776;
  assign T12776 = T12793 ? T12784 : twiddle4_2_256_imag;
  assign twiddle4_2_256_imag = T12779 + T12777;
  assign T12777 = $signed(T12778) / $signed(22'h100000);
  assign T12778 = $signed(32'h40000000) * $signed(16'hffff);
  assign T12779 = {T12782, T12780};
  assign T12780 = $signed(T12781) / $signed(22'h100000);
  assign T12781 = $signed(1'h0) * $signed(16'h0);
  assign T12782 = T12783 ? 31'h7fffffff : 31'h0;
  assign T12783 = T12780[5'h10:5'h10];
  assign T12784 = {T12792, twiddle4_2_257_imag};
  assign twiddle4_2_257_imag = T12787 + T12785;
  assign T12785 = $signed(T12786) / $signed(22'h100000);
  assign T12786 = $signed(31'h3fffb10b) * $signed(16'hffff);
  assign T12787 = {T12790, T12788};
  assign T12788 = $signed(T12789) / $signed(22'h100000);
  assign T12789 = $signed(24'h9b783d) * $signed(16'h0);
  assign T12790 = T12791 ? 7'h7f : 7'h0;
  assign T12791 = T12788[6'h27:6'h27];
  assign T12792 = twiddle4_2_257_imag[6'h2e:6'h2e];
  assign T12793 = T10817[1'h0:1'h0];
  assign T12794 = {T12811, T12795};
  assign T12795 = T12810 ? twiddle4_2_259_imag : twiddle4_2_258_imag;
  assign twiddle4_2_258_imag = T12798 + T12796;
  assign T12796 = $signed(T12797) / $signed(22'h100000);
  assign T12797 = $signed(31'h3ffec42d) * $signed(16'hffff);
  assign T12798 = {T12801, T12799};
  assign T12799 = $signed(T12800) / $signed(22'h100000);
  assign T12800 = $signed(25'h136f171) * $signed(16'h0);
  assign T12801 = T12802 ? 6'h3f : 6'h0;
  assign T12802 = T12799[6'h28:6'h28];
  assign twiddle4_2_259_imag = T12805 + T12803;
  assign T12803 = $signed(T12804) / $signed(22'h100000);
  assign T12804 = $signed(31'h3ffd3968) * $signed(16'hffff);
  assign T12805 = {T12808, T12806};
  assign T12806 = $signed(T12807) / $signed(22'h100000);
  assign T12807 = $signed(26'h2d26c95) * $signed(16'h0);
  assign T12808 = T12809 ? 5'h1f : 5'h0;
  assign T12809 = T12806[6'h29:6'h29];
  assign T12810 = T10817[1'h0:1'h0];
  assign T12811 = T12795[6'h2e:6'h2e];
  assign T12812 = T10817[1'h1:1'h1];
  assign T12813 = {T12848, T12814};
  assign T12814 = T12847 ? T12831 : T12815;
  assign T12815 = T12830 ? twiddle4_2_261_imag : twiddle4_2_260_imag;
  assign twiddle4_2_260_imag = T12818 + T12816;
  assign T12816 = $signed(T12817) / $signed(22'h100000);
  assign T12817 = $signed(31'h3ffb10c1) * $signed(16'hffff);
  assign T12818 = {T12821, T12819};
  assign T12819 = $signed(T12820) / $signed(22'h100000);
  assign T12820 = $signed(26'h26deaa1) * $signed(16'h0);
  assign T12821 = T12822 ? 5'h1f : 5'h0;
  assign T12822 = T12819[6'h29:6'h29];
  assign twiddle4_2_261_imag = T12825 + T12823;
  assign T12823 = $signed(T12824) / $signed(22'h100000);
  assign T12824 = $signed(31'h3ff84a3b) * $signed(16'hffff);
  assign T12825 = {T12828, T12826};
  assign T12826 = $signed(T12827) / $signed(22'h100000);
  assign T12827 = $signed(26'h2096c8d) * $signed(16'h0);
  assign T12828 = T12829 ? 5'h1f : 5'h0;
  assign T12829 = T12826[6'h29:6'h29];
  assign T12830 = T10817[1'h0:1'h0];
  assign T12831 = T12846 ? twiddle4_2_263_imag : twiddle4_2_262_imag;
  assign twiddle4_2_262_imag = T12834 + T12832;
  assign T12832 = $signed(T12833) / $signed(22'h100000);
  assign T12833 = $signed(31'h3ff4e5df) * $signed(16'hffff);
  assign T12834 = {T12837, T12835};
  assign T12835 = $signed(T12836) / $signed(22'h100000);
  assign T12836 = $signed(27'h5a4f352) * $signed(16'h0);
  assign T12837 = T12838 ? 4'hf : 4'h0;
  assign T12838 = T12835[6'h2a:6'h2a];
  assign twiddle4_2_263_imag = T12841 + T12839;
  assign T12839 = $signed(T12840) / $signed(22'h100000);
  assign T12840 = $signed(31'h3ff0e3b5) * $signed(16'hffff);
  assign T12841 = {T12844, T12842};
  assign T12842 = $signed(T12843) / $signed(22'h100000);
  assign T12843 = $signed(27'h5407fe6) * $signed(16'h0);
  assign T12844 = T12845 ? 4'hf : 4'h0;
  assign T12845 = T12842[6'h2a:6'h2a];
  assign T12846 = T10817[1'h0:1'h0];
  assign T12847 = T10817[1'h1:1'h1];
  assign T12848 = T12814[6'h2e:6'h2e];
  assign T12849 = T10817[2'h2:2'h2];
  assign T12850 = {T12921, T12851};
  assign T12851 = T12920 ? T12886 : T12852;
  assign T12852 = T12885 ? T12869 : T12853;
  assign T12853 = T12868 ? twiddle4_2_265_imag : twiddle4_2_264_imag;
  assign twiddle4_2_264_imag = T12856 + T12854;
  assign T12854 = $signed(T12855) / $signed(22'h100000);
  assign T12855 = $signed(31'h3fec43c6) * $signed(16'hffff);
  assign T12856 = {T12859, T12857};
  assign T12857 = $signed(T12858) / $signed(22'h100000);
  assign T12858 = $signed(27'h4dc1342) * $signed(16'h0);
  assign T12859 = T12860 ? 4'hf : 4'h0;
  assign T12860 = T12857[6'h2a:6'h2a];
  assign twiddle4_2_265_imag = T12863 + T12861;
  assign T12861 = $signed(T12862) / $signed(22'h100000);
  assign T12862 = $signed(31'h3fe7061f) * $signed(16'hffff);
  assign T12863 = {T12866, T12864};
  assign T12864 = $signed(T12865) / $signed(22'h100000);
  assign T12865 = $signed(27'h477ae5e) * $signed(16'h0);
  assign T12866 = T12867 ? 4'hf : 4'h0;
  assign T12867 = T12864[6'h2a:6'h2a];
  assign T12868 = T10817[1'h0:1'h0];
  assign T12869 = T12884 ? twiddle4_2_267_imag : twiddle4_2_266_imag;
  assign twiddle4_2_266_imag = T12872 + T12870;
  assign T12870 = $signed(T12871) / $signed(22'h100000);
  assign T12871 = $signed(31'h3fe12acb) * $signed(16'hffff);
  assign T12872 = {T12875, T12873};
  assign T12873 = $signed(T12874) / $signed(22'h100000);
  assign T12874 = $signed(27'h4135231) * $signed(16'h0);
  assign T12875 = T12876 ? 4'hf : 4'h0;
  assign T12876 = T12873[6'h2a:6'h2a];
  assign twiddle4_2_267_imag = T12879 + T12877;
  assign T12877 = $signed(T12878) / $signed(22'h100000);
  assign T12878 = $signed(31'h3fdab1d9) * $signed(16'hffff);
  assign T12879 = {T12882, T12880};
  assign T12880 = $signed(T12881) / $signed(22'h100000);
  assign T12881 = $signed(28'hbaeffb3) * $signed(16'h0);
  assign T12882 = T12883 ? 3'h7 : 3'h0;
  assign T12883 = T12880[6'h2b:6'h2b];
  assign T12884 = T10817[1'h0:1'h0];
  assign T12885 = T10817[1'h1:1'h1];
  assign T12886 = T12919 ? T12903 : T12887;
  assign T12887 = T12902 ? twiddle4_2_269_imag : twiddle4_2_268_imag;
  assign twiddle4_2_268_imag = T12890 + T12888;
  assign T12888 = $signed(T12889) / $signed(22'h100000);
  assign T12889 = $signed(31'h3fd39b5a) * $signed(16'hffff);
  assign T12890 = {T12893, T12891};
  assign T12891 = $signed(T12892) / $signed(22'h100000);
  assign T12892 = $signed(28'hb4ab7dc) * $signed(16'h0);
  assign T12893 = T12894 ? 3'h7 : 3'h0;
  assign T12894 = T12891[6'h2b:6'h2b];
  assign twiddle4_2_269_imag = T12897 + T12895;
  assign T12895 = $signed(T12896) / $signed(22'h100000);
  assign T12896 = $signed(31'h3fcbe75e) * $signed(16'hffff);
  assign T12897 = {T12900, T12898};
  assign T12898 = $signed(T12899) / $signed(22'h100000);
  assign T12899 = $signed(28'hae67ba2) * $signed(16'h0);
  assign T12900 = T12901 ? 3'h7 : 3'h0;
  assign T12901 = T12898[6'h2b:6'h2b];
  assign T12902 = T10817[1'h0:1'h0];
  assign T12903 = T12918 ? twiddle4_2_271_imag : twiddle4_2_270_imag;
  assign twiddle4_2_270_imag = T12906 + T12904;
  assign T12904 = $signed(T12905) / $signed(22'h100000);
  assign T12905 = $signed(31'h3fc395f9) * $signed(16'hffff);
  assign T12906 = {T12909, T12907};
  assign T12907 = $signed(T12908) / $signed(22'h100000);
  assign T12908 = $signed(28'ha824bfe) * $signed(16'h0);
  assign T12909 = T12910 ? 3'h7 : 3'h0;
  assign T12910 = T12907[6'h2b:6'h2b];
  assign twiddle4_2_271_imag = T12913 + T12911;
  assign T12911 = $signed(T12912) / $signed(22'h100000);
  assign T12912 = $signed(31'h3fbaa73f) * $signed(16'hffff);
  assign T12913 = {T12916, T12914};
  assign T12914 = $signed(T12915) / $signed(22'h100000);
  assign T12915 = $signed(28'ha1e29e6) * $signed(16'h0);
  assign T12916 = T12917 ? 3'h7 : 3'h0;
  assign T12917 = T12914[6'h2b:6'h2b];
  assign T12918 = T10817[1'h0:1'h0];
  assign T12919 = T10817[1'h1:1'h1];
  assign T12920 = T10817[2'h2:2'h2];
  assign T12921 = T12851[6'h2e:6'h2e];
  assign T12922 = T10817[2'h3:2'h3];
  assign T12923 = {T13066, T12924};
  assign T12924 = T13065 ? T12995 : T12925;
  assign T12925 = T12994 ? T12960 : T12926;
  assign T12926 = T12959 ? T12943 : T12927;
  assign T12927 = T12942 ? twiddle4_2_273_imag : twiddle4_2_272_imag;
  assign twiddle4_2_272_imag = T12930 + T12928;
  assign T12928 = $signed(T12929) / $signed(22'h100000);
  assign T12929 = $signed(31'h3fb11b47) * $signed(16'hffff);
  assign T12930 = {T12933, T12931};
  assign T12931 = $signed(T12932) / $signed(22'h100000);
  assign T12932 = $signed(28'h9ba1651) * $signed(16'h0);
  assign T12933 = T12934 ? 3'h7 : 3'h0;
  assign T12934 = T12931[6'h2b:6'h2b];
  assign twiddle4_2_273_imag = T12937 + T12935;
  assign T12935 = $signed(T12936) / $signed(22'h100000);
  assign T12936 = $signed(31'h3fa6f228) * $signed(16'hffff);
  assign T12937 = {T12940, T12938};
  assign T12938 = $signed(T12939) / $signed(22'h100000);
  assign T12939 = $signed(28'h9561237) * $signed(16'h0);
  assign T12940 = T12941 ? 3'h7 : 3'h0;
  assign T12941 = T12938[6'h2b:6'h2b];
  assign T12942 = T10817[1'h0:1'h0];
  assign T12943 = T12958 ? twiddle4_2_275_imag : twiddle4_2_274_imag;
  assign twiddle4_2_274_imag = T12946 + T12944;
  assign T12944 = $signed(T12945) / $signed(22'h100000);
  assign T12945 = $signed(31'h3f9c2bfa) * $signed(16'hffff);
  assign T12946 = {T12949, T12947};
  assign T12947 = $signed(T12948) / $signed(22'h100000);
  assign T12948 = $signed(28'h8f21e8f) * $signed(16'h0);
  assign T12949 = T12950 ? 3'h7 : 3'h0;
  assign T12950 = T12947[6'h2b:6'h2b];
  assign twiddle4_2_275_imag = T12953 + T12951;
  assign T12951 = $signed(T12952) / $signed(22'h100000);
  assign T12952 = $signed(31'h3f90c8d9) * $signed(16'hffff);
  assign T12953 = {T12956, T12954};
  assign T12954 = $signed(T12955) / $signed(22'h100000);
  assign T12955 = $signed(28'h88e3c4e) * $signed(16'h0);
  assign T12956 = T12957 ? 3'h7 : 3'h0;
  assign T12957 = T12954[6'h2b:6'h2b];
  assign T12958 = T10817[1'h0:1'h0];
  assign T12959 = T10817[1'h1:1'h1];
  assign T12960 = T12993 ? T12977 : T12961;
  assign T12961 = T12976 ? twiddle4_2_277_imag : twiddle4_2_276_imag;
  assign twiddle4_2_276_imag = T12964 + T12962;
  assign T12962 = $signed(T12963) / $signed(22'h100000);
  assign T12963 = $signed(31'h3f84c8e1) * $signed(16'hffff);
  assign T12964 = {T12967, T12965};
  assign T12965 = $signed(T12966) / $signed(22'h100000);
  assign T12966 = $signed(28'h82a6c6b) * $signed(16'h0);
  assign T12967 = T12968 ? 3'h7 : 3'h0;
  assign T12968 = T12965[6'h2b:6'h2b];
  assign twiddle4_2_277_imag = T12971 + T12969;
  assign T12969 = $signed(T12970) / $signed(22'h100000);
  assign T12970 = $signed(31'h3f782c2f) * $signed(16'hffff);
  assign T12971 = {T12974, T12972};
  assign T12972 = $signed(T12973) / $signed(22'h100000);
  assign T12973 = $signed(29'h17c6afdd) * $signed(16'h0);
  assign T12974 = T12975 ? 2'h3 : 2'h0;
  assign T12975 = T12972[6'h2c:6'h2c];
  assign T12976 = T10817[1'h0:1'h0];
  assign T12977 = T12992 ? twiddle4_2_279_imag : twiddle4_2_278_imag;
  assign twiddle4_2_278_imag = T12980 + T12978;
  assign T12978 = $signed(T12979) / $signed(22'h100000);
  assign T12979 = $signed(31'h3f6af2e3) * $signed(16'hffff);
  assign T12980 = {T12983, T12981};
  assign T12981 = $signed(T12982) / $signed(22'h100000);
  assign T12982 = $signed(29'h17630799) * $signed(16'h0);
  assign T12983 = T12984 ? 2'h3 : 2'h0;
  assign T12984 = T12981[6'h2c:6'h2c];
  assign twiddle4_2_279_imag = T12987 + T12985;
  assign T12985 = $signed(T12986) / $signed(22'h100000);
  assign T12986 = $signed(31'h3f5d1d1c) * $signed(16'hffff);
  assign T12987 = {T12990, T12988};
  assign T12988 = $signed(T12989) / $signed(22'h100000);
  assign T12989 = $signed(29'h16ff7496) * $signed(16'h0);
  assign T12990 = T12991 ? 2'h3 : 2'h0;
  assign T12991 = T12988[6'h2c:6'h2c];
  assign T12992 = T10817[1'h0:1'h0];
  assign T12993 = T10817[1'h1:1'h1];
  assign T12994 = T10817[2'h2:2'h2];
  assign T12995 = T13064 ? T13030 : T12996;
  assign T12996 = T13029 ? T13013 : T12997;
  assign T12997 = T13012 ? twiddle4_2_281_imag : twiddle4_2_280_imag;
  assign twiddle4_2_280_imag = T13000 + T12998;
  assign T12998 = $signed(T12999) / $signed(22'h100000);
  assign T12999 = $signed(31'h3f4eaafe) * $signed(16'hffff);
  assign T13000 = {T13003, T13001};
  assign T13001 = $signed(T13002) / $signed(22'h100000);
  assign T13002 = $signed(29'h169bf7c9) * $signed(16'h0);
  assign T13003 = T13004 ? 2'h3 : 2'h0;
  assign T13004 = T13001[6'h2c:6'h2c];
  assign twiddle4_2_281_imag = T13007 + T13005;
  assign T13005 = $signed(T13006) / $signed(22'h100000);
  assign T13006 = $signed(31'h3f3f9cab) * $signed(16'hffff);
  assign T13007 = {T13010, T13008};
  assign T13008 = $signed(T13009) / $signed(22'h100000);
  assign T13009 = $signed(29'h16389228) * $signed(16'h0);
  assign T13010 = T13011 ? 2'h3 : 2'h0;
  assign T13011 = T13008[6'h2c:6'h2c];
  assign T13012 = T10817[1'h0:1'h0];
  assign T13013 = T13028 ? twiddle4_2_283_imag : twiddle4_2_282_imag;
  assign twiddle4_2_282_imag = T13016 + T13014;
  assign T13014 = $signed(T13015) / $signed(22'h100000);
  assign T13015 = $signed(31'h3f2ff249) * $signed(16'hffff);
  assign T13016 = {T13019, T13017};
  assign T13017 = $signed(T13018) / $signed(22'h100000);
  assign T13018 = $signed(29'h15d544a8) * $signed(16'h0);
  assign T13019 = T13020 ? 2'h3 : 2'h0;
  assign T13020 = T13017[6'h2c:6'h2c];
  assign twiddle4_2_283_imag = T13023 + T13021;
  assign T13021 = $signed(T13022) / $signed(22'h100000);
  assign T13022 = $signed(31'h3f1fabff) * $signed(16'hffff);
  assign T13023 = {T13026, T13024};
  assign T13024 = $signed(T13025) / $signed(22'h100000);
  assign T13025 = $signed(29'h1572103e) * $signed(16'h0);
  assign T13026 = T13027 ? 2'h3 : 2'h0;
  assign T13027 = T13024[6'h2c:6'h2c];
  assign T13028 = T10817[1'h0:1'h0];
  assign T13029 = T10817[1'h1:1'h1];
  assign T13030 = T13063 ? T13047 : T13031;
  assign T13031 = T13046 ? twiddle4_2_285_imag : twiddle4_2_284_imag;
  assign twiddle4_2_284_imag = T13034 + T13032;
  assign T13032 = $signed(T13033) / $signed(22'h100000);
  assign T13033 = $signed(31'h3f0ec9f4) * $signed(16'hffff);
  assign T13034 = {T13037, T13035};
  assign T13035 = $signed(T13036) / $signed(22'h100000);
  assign T13036 = $signed(29'h150ef5de) * $signed(16'h0);
  assign T13037 = T13038 ? 2'h3 : 2'h0;
  assign T13038 = T13035[6'h2c:6'h2c];
  assign twiddle4_2_285_imag = T13041 + T13039;
  assign T13039 = $signed(T13040) / $signed(22'h100000);
  assign T13040 = $signed(31'h3efd4c53) * $signed(16'hffff);
  assign T13041 = {T13044, T13042};
  assign T13042 = $signed(T13043) / $signed(22'h100000);
  assign T13043 = $signed(29'h14abf67e) * $signed(16'h0);
  assign T13044 = T13045 ? 2'h3 : 2'h0;
  assign T13045 = T13042[6'h2c:6'h2c];
  assign T13046 = T10817[1'h0:1'h0];
  assign T13047 = T13062 ? twiddle4_2_287_imag : twiddle4_2_286_imag;
  assign twiddle4_2_286_imag = T13050 + T13048;
  assign T13048 = $signed(T13049) / $signed(22'h100000);
  assign T13049 = $signed(31'h3eeb3347) * $signed(16'hffff);
  assign T13050 = {T13053, T13051};
  assign T13051 = $signed(T13052) / $signed(22'h100000);
  assign T13052 = $signed(29'h14491311) * $signed(16'h0);
  assign T13053 = T13054 ? 2'h3 : 2'h0;
  assign T13054 = T13051[6'h2c:6'h2c];
  assign twiddle4_2_287_imag = T13057 + T13055;
  assign T13055 = $signed(T13056) / $signed(22'h100000);
  assign T13056 = $signed(31'h3ed87efb) * $signed(16'hffff);
  assign T13057 = {T13060, T13058};
  assign T13058 = $signed(T13059) / $signed(22'h100000);
  assign T13059 = $signed(29'h13e64c8c) * $signed(16'h0);
  assign T13060 = T13061 ? 2'h3 : 2'h0;
  assign T13061 = T13058[6'h2c:6'h2c];
  assign T13062 = T10817[1'h0:1'h0];
  assign T13063 = T10817[1'h1:1'h1];
  assign T13064 = T10817[2'h2:2'h2];
  assign T13065 = T10817[2'h3:2'h3];
  assign T13066 = T12924[6'h2e:6'h2e];
  assign T13067 = T10817[3'h4:3'h4];
  assign T13068 = {T13333, T13069};
  assign T13069 = T13332 ? T13206 : T13070;
  assign T13070 = T13205 ? T13141 : T13071;
  assign T13071 = T13140 ? T13106 : T13072;
  assign T13072 = T13105 ? T13089 : T13073;
  assign T13073 = T13088 ? twiddle4_2_289_imag : twiddle4_2_288_imag;
  assign twiddle4_2_288_imag = T13076 + T13074;
  assign T13074 = $signed(T13075) / $signed(22'h100000);
  assign T13075 = $signed(31'h3ec52f9f) * $signed(16'hffff);
  assign T13076 = {T13079, T13077};
  assign T13077 = $signed(T13078) / $signed(22'h100000);
  assign T13078 = $signed(29'h1383a3e2) * $signed(16'h0);
  assign T13079 = T13080 ? 2'h3 : 2'h0;
  assign T13080 = T13077[6'h2c:6'h2c];
  assign twiddle4_2_289_imag = T13083 + T13081;
  assign T13081 = $signed(T13082) / $signed(22'h100000);
  assign T13082 = $signed(31'h3eb14562) * $signed(16'hffff);
  assign T13083 = {T13086, T13084};
  assign T13084 = $signed(T13085) / $signed(22'h100000);
  assign T13085 = $signed(29'h13211a07) * $signed(16'h0);
  assign T13086 = T13087 ? 2'h3 : 2'h0;
  assign T13087 = T13084[6'h2c:6'h2c];
  assign T13088 = T10817[1'h0:1'h0];
  assign T13089 = T13104 ? twiddle4_2_291_imag : twiddle4_2_290_imag;
  assign twiddle4_2_290_imag = T13092 + T13090;
  assign T13090 = $signed(T13091) / $signed(22'h100000);
  assign T13091 = $signed(31'h3e9cc076) * $signed(16'hffff);
  assign T13092 = {T13095, T13093};
  assign T13093 = $signed(T13094) / $signed(22'h100000);
  assign T13094 = $signed(29'h12beafee) * $signed(16'h0);
  assign T13095 = T13096 ? 2'h3 : 2'h0;
  assign T13096 = T13093[6'h2c:6'h2c];
  assign twiddle4_2_291_imag = T13099 + T13097;
  assign T13097 = $signed(T13098) / $signed(22'h100000);
  assign T13098 = $signed(31'h3e87a10b) * $signed(16'hffff);
  assign T13099 = {T13102, T13100};
  assign T13100 = $signed(T13101) / $signed(22'h100000);
  assign T13101 = $signed(29'h125c6689) * $signed(16'h0);
  assign T13102 = T13103 ? 2'h3 : 2'h0;
  assign T13103 = T13100[6'h2c:6'h2c];
  assign T13104 = T10817[1'h0:1'h0];
  assign T13105 = T10817[1'h1:1'h1];
  assign T13106 = T13139 ? T13123 : T13107;
  assign T13107 = T13122 ? twiddle4_2_293_imag : twiddle4_2_292_imag;
  assign twiddle4_2_292_imag = T13110 + T13108;
  assign T13108 = $signed(T13109) / $signed(22'h100000);
  assign T13109 = $signed(31'h3e71e758) * $signed(16'hffff);
  assign T13110 = {T13113, T13111};
  assign T13111 = $signed(T13112) / $signed(22'h100000);
  assign T13112 = $signed(29'h11fa3ecb) * $signed(16'h0);
  assign T13113 = T13114 ? 2'h3 : 2'h0;
  assign T13114 = T13111[6'h2c:6'h2c];
  assign twiddle4_2_293_imag = T13117 + T13115;
  assign T13115 = $signed(T13116) / $signed(22'h100000);
  assign T13116 = $signed(31'h3e5b9392) * $signed(16'hffff);
  assign T13117 = {T13120, T13118};
  assign T13118 = $signed(T13119) / $signed(22'h100000);
  assign T13119 = $signed(29'h119839a7) * $signed(16'h0);
  assign T13120 = T13121 ? 2'h3 : 2'h0;
  assign T13121 = T13118[6'h2c:6'h2c];
  assign T13122 = T10817[1'h0:1'h0];
  assign T13123 = T13138 ? twiddle4_2_295_imag : twiddle4_2_294_imag;
  assign twiddle4_2_294_imag = T13126 + T13124;
  assign T13124 = $signed(T13125) / $signed(22'h100000);
  assign T13125 = $signed(31'h3e44a5ee) * $signed(16'hffff);
  assign T13126 = {T13129, T13127};
  assign T13127 = $signed(T13128) / $signed(22'h100000);
  assign T13128 = $signed(29'h1136580e) * $signed(16'h0);
  assign T13129 = T13130 ? 2'h3 : 2'h0;
  assign T13130 = T13127[6'h2c:6'h2c];
  assign twiddle4_2_295_imag = T13133 + T13131;
  assign T13131 = $signed(T13132) / $signed(22'h100000);
  assign T13132 = $signed(31'h3e2d1ea7) * $signed(16'hffff);
  assign T13133 = {T13136, T13134};
  assign T13134 = $signed(T13135) / $signed(22'h100000);
  assign T13135 = $signed(29'h10d49af1) * $signed(16'h0);
  assign T13136 = T13137 ? 2'h3 : 2'h0;
  assign T13137 = T13134[6'h2c:6'h2c];
  assign T13138 = T10817[1'h0:1'h0];
  assign T13139 = T10817[1'h1:1'h1];
  assign T13140 = T10817[2'h2:2'h2];
  assign T13141 = T13204 ? T13174 : T13142;
  assign T13142 = T13173 ? T13159 : T13143;
  assign T13143 = T13158 ? twiddle4_2_297_imag : twiddle4_2_296_imag;
  assign twiddle4_2_296_imag = T13146 + T13144;
  assign T13144 = $signed(T13145) / $signed(22'h100000);
  assign T13145 = $signed(31'h3e14fdf7) * $signed(16'hffff);
  assign T13146 = {T13149, T13147};
  assign T13147 = $signed(T13148) / $signed(22'h100000);
  assign T13148 = $signed(29'h10730343) * $signed(16'h0);
  assign T13149 = T13150 ? 2'h3 : 2'h0;
  assign T13150 = T13147[6'h2c:6'h2c];
  assign twiddle4_2_297_imag = T13153 + T13151;
  assign T13151 = $signed(T13152) / $signed(22'h100000);
  assign T13152 = $signed(31'h3dfc4418) * $signed(16'hffff);
  assign T13153 = {T13156, T13154};
  assign T13154 = $signed(T13155) / $signed(22'h100000);
  assign T13155 = $signed(29'h101191f3) * $signed(16'h0);
  assign T13156 = T13157 ? 2'h3 : 2'h0;
  assign T13157 = T13154[6'h2c:6'h2c];
  assign T13158 = T10817[1'h0:1'h0];
  assign T13159 = T13172 ? twiddle4_2_299_imag : twiddle4_2_298_imag;
  assign twiddle4_2_298_imag = T13162 + T13160;
  assign T13160 = $signed(T13161) / $signed(22'h100000);
  assign T13161 = $signed(31'h3de2f147) * $signed(16'hffff);
  assign T13162 = {T13165, T13163};
  assign T13163 = $signed(T13164) / $signed(22'h100000);
  assign T13164 = $signed(30'h2fb047f2) * $signed(16'h0);
  assign T13165 = T13163[6'h2d:6'h2d];
  assign twiddle4_2_299_imag = T13168 + T13166;
  assign T13166 = $signed(T13167) / $signed(22'h100000);
  assign T13167 = $signed(31'h3dc905c4) * $signed(16'hffff);
  assign T13168 = {T13171, T13169};
  assign T13169 = $signed(T13170) / $signed(22'h100000);
  assign T13170 = $signed(30'h2f4f2631) * $signed(16'h0);
  assign T13171 = T13169[6'h2d:6'h2d];
  assign T13172 = T10817[1'h0:1'h0];
  assign T13173 = T10817[1'h1:1'h1];
  assign T13174 = T13203 ? T13189 : T13175;
  assign T13175 = T13188 ? twiddle4_2_301_imag : twiddle4_2_300_imag;
  assign twiddle4_2_300_imag = T13178 + T13176;
  assign T13176 = $signed(T13177) / $signed(22'h100000);
  assign T13177 = $signed(31'h3dae81ce) * $signed(16'hffff);
  assign T13178 = {T13181, T13179};
  assign T13179 = $signed(T13180) / $signed(22'h100000);
  assign T13180 = $signed(30'h2eee2d9e) * $signed(16'h0);
  assign T13181 = T13179[6'h2d:6'h2d];
  assign twiddle4_2_301_imag = T13184 + T13182;
  assign T13182 = $signed(T13183) / $signed(22'h100000);
  assign T13183 = $signed(31'h3d9365a7) * $signed(16'hffff);
  assign T13184 = {T13187, T13185};
  assign T13185 = $signed(T13186) / $signed(22'h100000);
  assign T13186 = $signed(30'h2e8d5f29) * $signed(16'h0);
  assign T13187 = T13185[6'h2d:6'h2d];
  assign T13188 = T10817[1'h0:1'h0];
  assign T13189 = T13202 ? twiddle4_2_303_imag : twiddle4_2_302_imag;
  assign twiddle4_2_302_imag = T13192 + T13190;
  assign T13190 = $signed(T13191) / $signed(22'h100000);
  assign T13191 = $signed(31'h3d77b191) * $signed(16'hffff);
  assign T13192 = {T13195, T13193};
  assign T13193 = $signed(T13194) / $signed(22'h100000);
  assign T13194 = $signed(30'h2e2cbbc1) * $signed(16'h0);
  assign T13195 = T13193[6'h2d:6'h2d];
  assign twiddle4_2_303_imag = T13198 + T13196;
  assign T13196 = $signed(T13197) / $signed(22'h100000);
  assign T13197 = $signed(31'h3d5b65d1) * $signed(16'hffff);
  assign T13198 = {T13201, T13199};
  assign T13199 = $signed(T13200) / $signed(22'h100000);
  assign T13200 = $signed(30'h2dcc4455) * $signed(16'h0);
  assign T13201 = T13199[6'h2d:6'h2d];
  assign T13202 = T10817[1'h0:1'h0];
  assign T13203 = T10817[1'h1:1'h1];
  assign T13204 = T10817[2'h2:2'h2];
  assign T13205 = T10817[2'h3:2'h3];
  assign T13206 = T13331 ? T13269 : T13207;
  assign T13207 = T13268 ? T13238 : T13208;
  assign T13208 = T13237 ? T13223 : T13209;
  assign T13209 = T13222 ? twiddle4_2_305_imag : twiddle4_2_304_imag;
  assign twiddle4_2_304_imag = T13212 + T13210;
  assign T13210 = $signed(T13211) / $signed(22'h100000);
  assign T13211 = $signed(31'h3d3e82ad) * $signed(16'hffff);
  assign T13212 = {T13215, T13213};
  assign T13213 = $signed(T13214) / $signed(22'h100000);
  assign T13214 = $signed(30'h2d6bf9d2) * $signed(16'h0);
  assign T13215 = T13213[6'h2d:6'h2d];
  assign twiddle4_2_305_imag = T13218 + T13216;
  assign T13216 = $signed(T13217) / $signed(22'h100000);
  assign T13217 = $signed(31'h3d21086c) * $signed(16'hffff);
  assign T13218 = {T13221, T13219};
  assign T13219 = $signed(T13220) / $signed(22'h100000);
  assign T13220 = $signed(30'h2d0bdd26) * $signed(16'h0);
  assign T13221 = T13219[6'h2d:6'h2d];
  assign T13222 = T10817[1'h0:1'h0];
  assign T13223 = T13236 ? twiddle4_2_307_imag : twiddle4_2_306_imag;
  assign twiddle4_2_306_imag = T13226 + T13224;
  assign T13224 = $signed(T13225) / $signed(22'h100000);
  assign T13225 = $signed(31'h3d02f756) * $signed(16'hffff);
  assign T13226 = {T13229, T13227};
  assign T13227 = $signed(T13228) / $signed(22'h100000);
  assign T13228 = $signed(30'h2cabef3e) * $signed(16'h0);
  assign T13229 = T13227[6'h2d:6'h2d];
  assign twiddle4_2_307_imag = T13232 + T13230;
  assign T13230 = $signed(T13231) / $signed(22'h100000);
  assign T13231 = $signed(31'h3ce44fb6) * $signed(16'hffff);
  assign T13232 = {T13235, T13233};
  assign T13233 = $signed(T13234) / $signed(22'h100000);
  assign T13234 = $signed(30'h2c4c3106) * $signed(16'h0);
  assign T13235 = T13233[6'h2d:6'h2d];
  assign T13236 = T10817[1'h0:1'h0];
  assign T13237 = T10817[1'h1:1'h1];
  assign T13238 = T13267 ? T13253 : T13239;
  assign T13239 = T13252 ? twiddle4_2_309_imag : twiddle4_2_308_imag;
  assign twiddle4_2_308_imag = T13242 + T13240;
  assign T13240 = $signed(T13241) / $signed(22'h100000);
  assign T13241 = $signed(31'h3cc511d8) * $signed(16'hffff);
  assign T13242 = {T13245, T13243};
  assign T13243 = $signed(T13244) / $signed(22'h100000);
  assign T13244 = $signed(30'h2beca36c) * $signed(16'h0);
  assign T13245 = T13243[6'h2d:6'h2d];
  assign twiddle4_2_309_imag = T13248 + T13246;
  assign T13246 = $signed(T13247) / $signed(22'h100000);
  assign T13247 = $signed(31'h3ca53e08) * $signed(16'hffff);
  assign T13248 = {T13251, T13249};
  assign T13249 = $signed(T13250) / $signed(22'h100000);
  assign T13250 = $signed(30'h2b8d475b) * $signed(16'h0);
  assign T13251 = T13249[6'h2d:6'h2d];
  assign T13252 = T10817[1'h0:1'h0];
  assign T13253 = T13266 ? twiddle4_2_311_imag : twiddle4_2_310_imag;
  assign twiddle4_2_310_imag = T13256 + T13254;
  assign T13254 = $signed(T13255) / $signed(22'h100000);
  assign T13255 = $signed(31'h3c84d496) * $signed(16'hffff);
  assign T13256 = {T13259, T13257};
  assign T13257 = $signed(T13258) / $signed(22'h100000);
  assign T13258 = $signed(30'h2b2e1dbe) * $signed(16'h0);
  assign T13259 = T13257[6'h2d:6'h2d];
  assign twiddle4_2_311_imag = T13262 + T13260;
  assign T13260 = $signed(T13261) / $signed(22'h100000);
  assign T13261 = $signed(31'h3c63d5d0) * $signed(16'hffff);
  assign T13262 = {T13265, T13263};
  assign T13263 = $signed(T13264) / $signed(22'h100000);
  assign T13264 = $signed(30'h2acf2780) * $signed(16'h0);
  assign T13265 = T13263[6'h2d:6'h2d];
  assign T13266 = T10817[1'h0:1'h0];
  assign T13267 = T10817[1'h1:1'h1];
  assign T13268 = T10817[2'h2:2'h2];
  assign T13269 = T13330 ? T13300 : T13270;
  assign T13270 = T13299 ? T13285 : T13271;
  assign T13271 = T13284 ? twiddle4_2_313_imag : twiddle4_2_312_imag;
  assign twiddle4_2_312_imag = T13274 + T13272;
  assign T13272 = $signed(T13273) / $signed(22'h100000);
  assign T13273 = $signed(31'h3c424209) * $signed(16'hffff);
  assign T13274 = {T13277, T13275};
  assign T13275 = $signed(T13276) / $signed(22'h100000);
  assign T13276 = $signed(30'h2a70658b) * $signed(16'h0);
  assign T13277 = T13275[6'h2d:6'h2d];
  assign twiddle4_2_313_imag = T13280 + T13278;
  assign T13278 = $signed(T13279) / $signed(22'h100000);
  assign T13279 = $signed(31'h3c201994) * $signed(16'hffff);
  assign T13280 = {T13283, T13281};
  assign T13281 = $signed(T13282) / $signed(22'h100000);
  assign T13282 = $signed(30'h2a11d8c9) * $signed(16'h0);
  assign T13283 = T13281[6'h2d:6'h2d];
  assign T13284 = T10817[1'h0:1'h0];
  assign T13285 = T13298 ? twiddle4_2_315_imag : twiddle4_2_314_imag;
  assign twiddle4_2_314_imag = T13288 + T13286;
  assign T13286 = $signed(T13287) / $signed(22'h100000);
  assign T13287 = $signed(31'h3bfd5cc4) * $signed(16'hffff);
  assign T13288 = {T13291, T13289};
  assign T13289 = $signed(T13290) / $signed(22'h100000);
  assign T13290 = $signed(30'h29b38223) * $signed(16'h0);
  assign T13291 = T13289[6'h2d:6'h2d];
  assign twiddle4_2_315_imag = T13294 + T13292;
  assign T13292 = $signed(T13293) / $signed(22'h100000);
  assign T13293 = $signed(31'h3bda0bef) * $signed(16'hffff);
  assign T13294 = {T13297, T13295};
  assign T13295 = $signed(T13296) / $signed(22'h100000);
  assign T13296 = $signed(30'h29556283) * $signed(16'h0);
  assign T13297 = T13295[6'h2d:6'h2d];
  assign T13298 = T10817[1'h0:1'h0];
  assign T13299 = T10817[1'h1:1'h1];
  assign T13300 = T13329 ? T13315 : T13301;
  assign T13301 = T13314 ? twiddle4_2_317_imag : twiddle4_2_316_imag;
  assign twiddle4_2_316_imag = T13304 + T13302;
  assign T13302 = $signed(T13303) / $signed(22'h100000);
  assign T13303 = $signed(31'h3bb6276d) * $signed(16'hffff);
  assign T13304 = {T13307, T13305};
  assign T13305 = $signed(T13306) / $signed(22'h100000);
  assign T13306 = $signed(30'h28f77ad0) * $signed(16'h0);
  assign T13307 = T13305[6'h2d:6'h2d];
  assign twiddle4_2_317_imag = T13310 + T13308;
  assign T13308 = $signed(T13309) / $signed(22'h100000);
  assign T13309 = $signed(31'h3b91af96) * $signed(16'hffff);
  assign T13310 = {T13313, T13311};
  assign T13311 = $signed(T13312) / $signed(22'h100000);
  assign T13312 = $signed(30'h2899cbf1) * $signed(16'h0);
  assign T13313 = T13311[6'h2d:6'h2d];
  assign T13314 = T10817[1'h0:1'h0];
  assign T13315 = T13328 ? twiddle4_2_319_imag : twiddle4_2_318_imag;
  assign twiddle4_2_318_imag = T13318 + T13316;
  assign T13316 = $signed(T13317) / $signed(22'h100000);
  assign T13317 = $signed(31'h3b6ca4c4) * $signed(16'hffff);
  assign T13318 = {T13321, T13319};
  assign T13319 = $signed(T13320) / $signed(22'h100000);
  assign T13320 = $signed(30'h283c56cf) * $signed(16'h0);
  assign T13321 = T13319[6'h2d:6'h2d];
  assign twiddle4_2_319_imag = T13324 + T13322;
  assign T13322 = $signed(T13323) / $signed(22'h100000);
  assign T13323 = $signed(31'h3b470752) * $signed(16'hffff);
  assign T13324 = {T13327, T13325};
  assign T13325 = $signed(T13326) / $signed(22'h100000);
  assign T13326 = $signed(30'h27df1c50) * $signed(16'h0);
  assign T13327 = T13325[6'h2d:6'h2d];
  assign T13328 = T10817[1'h0:1'h0];
  assign T13329 = T10817[1'h1:1'h1];
  assign T13330 = T10817[2'h2:2'h2];
  assign T13331 = T10817[2'h3:2'h3];
  assign T13332 = T10817[3'h4:3'h4];
  assign T13333 = T13069[6'h2e:6'h2e];
  assign T13334 = T10817[3'h5:3'h5];
  assign T13335 = {T13762, T13336};
  assign T13336 = T13761 ? T13571 : T13337;
  assign T13337 = T13570 ? T13464 : T13338;
  assign T13338 = T13463 ? T13401 : T13339;
  assign T13339 = T13400 ? T13370 : T13340;
  assign T13340 = T13369 ? T13355 : T13341;
  assign T13341 = T13354 ? twiddle4_2_321_imag : twiddle4_2_320_imag;
  assign twiddle4_2_320_imag = T13344 + T13342;
  assign T13342 = $signed(T13343) / $signed(22'h100000);
  assign T13343 = $signed(31'h3b20d79e) * $signed(16'hffff);
  assign T13344 = {T13347, T13345};
  assign T13345 = $signed(T13346) / $signed(22'h100000);
  assign T13346 = $signed(30'h27821d5a) * $signed(16'h0);
  assign T13347 = T13345[6'h2d:6'h2d];
  assign twiddle4_2_321_imag = T13350 + T13348;
  assign T13348 = $signed(T13349) / $signed(22'h100000);
  assign T13349 = $signed(31'h3afa1605) * $signed(16'hffff);
  assign T13350 = {T13353, T13351};
  assign T13351 = $signed(T13352) / $signed(22'h100000);
  assign T13352 = $signed(30'h27255ad2) * $signed(16'h0);
  assign T13353 = T13351[6'h2d:6'h2d];
  assign T13354 = T10817[1'h0:1'h0];
  assign T13355 = T13368 ? twiddle4_2_323_imag : twiddle4_2_322_imag;
  assign twiddle4_2_322_imag = T13358 + T13356;
  assign T13356 = $signed(T13357) / $signed(22'h100000);
  assign T13357 = $signed(31'h3ad2c2e7) * $signed(16'hffff);
  assign T13358 = {T13361, T13359};
  assign T13359 = $signed(T13360) / $signed(22'h100000);
  assign T13360 = $signed(30'h26c8d59d) * $signed(16'h0);
  assign T13361 = T13359[6'h2d:6'h2d];
  assign twiddle4_2_323_imag = T13364 + T13362;
  assign T13362 = $signed(T13363) / $signed(22'h100000);
  assign T13363 = $signed(31'h3aaadea5) * $signed(16'hffff);
  assign T13364 = {T13367, T13365};
  assign T13365 = $signed(T13366) / $signed(22'h100000);
  assign T13366 = $signed(30'h266c8e9f) * $signed(16'h0);
  assign T13367 = T13365[6'h2d:6'h2d];
  assign T13368 = T10817[1'h0:1'h0];
  assign T13369 = T10817[1'h1:1'h1];
  assign T13370 = T13399 ? T13385 : T13371;
  assign T13371 = T13384 ? twiddle4_2_325_imag : twiddle4_2_324_imag;
  assign twiddle4_2_324_imag = T13374 + T13372;
  assign T13372 = $signed(T13373) / $signed(22'h100000);
  assign T13373 = $signed(31'h3a8269a2) * $signed(16'hffff);
  assign T13374 = {T13377, T13375};
  assign T13375 = $signed(T13376) / $signed(22'h100000);
  assign T13376 = $signed(30'h261086bd) * $signed(16'h0);
  assign T13377 = T13375[6'h2d:6'h2d];
  assign twiddle4_2_325_imag = T13380 + T13378;
  assign T13378 = $signed(T13379) / $signed(22'h100000);
  assign T13379 = $signed(31'h3a596441) * $signed(16'hffff);
  assign T13380 = {T13383, T13381};
  assign T13381 = $signed(T13382) / $signed(22'h100000);
  assign T13382 = $signed(30'h25b4bed9) * $signed(16'h0);
  assign T13383 = T13381[6'h2d:6'h2d];
  assign T13384 = T10817[1'h0:1'h0];
  assign T13385 = T13398 ? twiddle4_2_327_imag : twiddle4_2_326_imag;
  assign twiddle4_2_326_imag = T13388 + T13386;
  assign T13386 = $signed(T13387) / $signed(22'h100000);
  assign T13387 = $signed(31'h3a2fcee8) * $signed(16'hffff);
  assign T13388 = {T13391, T13389};
  assign T13389 = $signed(T13390) / $signed(22'h100000);
  assign T13390 = $signed(30'h255937d5) * $signed(16'h0);
  assign T13391 = T13389[6'h2d:6'h2d];
  assign twiddle4_2_327_imag = T13394 + T13392;
  assign T13392 = $signed(T13393) / $signed(22'h100000);
  assign T13393 = $signed(31'h3a05a9fd) * $signed(16'hffff);
  assign T13394 = {T13397, T13395};
  assign T13395 = $signed(T13396) / $signed(22'h100000);
  assign T13396 = $signed(30'h24fdf294) * $signed(16'h0);
  assign T13397 = T13395[6'h2d:6'h2d];
  assign T13398 = T10817[1'h0:1'h0];
  assign T13399 = T10817[1'h1:1'h1];
  assign T13400 = T10817[2'h2:2'h2];
  assign T13401 = T13462 ? T13432 : T13402;
  assign T13402 = T13431 ? T13417 : T13403;
  assign T13403 = T13416 ? twiddle4_2_329_imag : twiddle4_2_328_imag;
  assign twiddle4_2_328_imag = T13406 + T13404;
  assign T13404 = $signed(T13405) / $signed(22'h100000);
  assign T13405 = $signed(31'h39daf5e8) * $signed(16'hffff);
  assign T13406 = {T13409, T13407};
  assign T13407 = $signed(T13408) / $signed(22'h100000);
  assign T13408 = $signed(30'h24a2eff7) * $signed(16'h0);
  assign T13409 = T13407[6'h2d:6'h2d];
  assign twiddle4_2_329_imag = T13412 + T13410;
  assign T13410 = $signed(T13411) / $signed(22'h100000);
  assign T13411 = $signed(31'h39afb313) * $signed(16'hffff);
  assign T13412 = {T13415, T13413};
  assign T13413 = $signed(T13414) / $signed(22'h100000);
  assign T13414 = $signed(30'h244830dd) * $signed(16'h0);
  assign T13415 = T13413[6'h2d:6'h2d];
  assign T13416 = T10817[1'h0:1'h0];
  assign T13417 = T13430 ? twiddle4_2_331_imag : twiddle4_2_330_imag;
  assign twiddle4_2_330_imag = T13420 + T13418;
  assign T13418 = $signed(T13419) / $signed(22'h100000);
  assign T13419 = $signed(31'h3983e1e7) * $signed(16'hffff);
  assign T13420 = {T13423, T13421};
  assign T13421 = $signed(T13422) / $signed(22'h100000);
  assign T13422 = $signed(30'h23edb628) * $signed(16'h0);
  assign T13423 = T13421[6'h2d:6'h2d];
  assign twiddle4_2_331_imag = T13426 + T13424;
  assign T13424 = $signed(T13425) / $signed(22'h100000);
  assign T13425 = $signed(31'h395782d3) * $signed(16'hffff);
  assign T13426 = {T13429, T13427};
  assign T13427 = $signed(T13428) / $signed(22'h100000);
  assign T13428 = $signed(30'h239380b7) * $signed(16'h0);
  assign T13429 = T13427[6'h2d:6'h2d];
  assign T13430 = T10817[1'h0:1'h0];
  assign T13431 = T10817[1'h1:1'h1];
  assign T13432 = T13461 ? T13447 : T13433;
  assign T13433 = T13446 ? twiddle4_2_333_imag : twiddle4_2_332_imag;
  assign twiddle4_2_332_imag = T13436 + T13434;
  assign T13434 = $signed(T13435) / $signed(22'h100000);
  assign T13435 = $signed(31'h392a9642) * $signed(16'hffff);
  assign T13436 = {T13439, T13437};
  assign T13437 = $signed(T13438) / $signed(22'h100000);
  assign T13438 = $signed(30'h23399167) * $signed(16'h0);
  assign T13439 = T13437[6'h2d:6'h2d];
  assign twiddle4_2_333_imag = T13442 + T13440;
  assign T13440 = $signed(T13441) / $signed(22'h100000);
  assign T13441 = $signed(31'h38fd1ca4) * $signed(16'hffff);
  assign T13442 = {T13445, T13443};
  assign T13443 = $signed(T13444) / $signed(22'h100000);
  assign T13444 = $signed(30'h22dfe918) * $signed(16'h0);
  assign T13445 = T13443[6'h2d:6'h2d];
  assign T13446 = T10817[1'h0:1'h0];
  assign T13447 = T13460 ? twiddle4_2_335_imag : twiddle4_2_334_imag;
  assign twiddle4_2_334_imag = T13450 + T13448;
  assign T13448 = $signed(T13449) / $signed(22'h100000);
  assign T13449 = $signed(31'h38cf1669) * $signed(16'hffff);
  assign T13450 = {T13453, T13451};
  assign T13451 = $signed(T13452) / $signed(22'h100000);
  assign T13452 = $signed(30'h228688a5) * $signed(16'h0);
  assign T13453 = T13451[6'h2d:6'h2d];
  assign twiddle4_2_335_imag = T13456 + T13454;
  assign T13454 = $signed(T13455) / $signed(22'h100000);
  assign T13455 = $signed(31'h38a08402) * $signed(16'hffff);
  assign T13456 = {T13459, T13457};
  assign T13457 = $signed(T13458) / $signed(22'h100000);
  assign T13458 = $signed(30'h222d70ec) * $signed(16'h0);
  assign T13459 = T13457[6'h2d:6'h2d];
  assign T13460 = T10817[1'h0:1'h0];
  assign T13461 = T10817[1'h1:1'h1];
  assign T13462 = T10817[2'h2:2'h2];
  assign T13463 = T10817[2'h3:2'h3];
  assign T13464 = T13569 ? T13523 : T13465;
  assign T13465 = T13522 ? T13496 : T13466;
  assign T13466 = T13495 ? T13481 : T13467;
  assign T13467 = T13480 ? twiddle4_2_337_imag : twiddle4_2_336_imag;
  assign twiddle4_2_336_imag = T13470 + T13468;
  assign T13468 = $signed(T13469) / $signed(22'h100000);
  assign T13469 = $signed(31'h387165e3) * $signed(16'hffff);
  assign T13470 = {T13473, T13471};
  assign T13471 = $signed(T13472) / $signed(22'h100000);
  assign T13472 = $signed(30'h21d4a2c8) * $signed(16'h0);
  assign T13473 = T13471[6'h2d:6'h2d];
  assign twiddle4_2_337_imag = T13476 + T13474;
  assign T13474 = $signed(T13475) / $signed(22'h100000);
  assign T13475 = $signed(31'h3841bc7f) * $signed(16'hffff);
  assign T13476 = {T13479, T13477};
  assign T13477 = $signed(T13478) / $signed(22'h100000);
  assign T13478 = $signed(30'h217c1f16) * $signed(16'h0);
  assign T13479 = T13477[6'h2d:6'h2d];
  assign T13480 = T10817[1'h0:1'h0];
  assign T13481 = T13494 ? twiddle4_2_339_imag : twiddle4_2_338_imag;
  assign twiddle4_2_338_imag = T13484 + T13482;
  assign T13482 = $signed(T13483) / $signed(22'h100000);
  assign T13483 = $signed(31'h3811884c) * $signed(16'hffff);
  assign T13484 = {T13487, T13485};
  assign T13485 = $signed(T13486) / $signed(22'h100000);
  assign T13486 = $signed(30'h2123e6ae) * $signed(16'h0);
  assign T13487 = T13485[6'h2d:6'h2d];
  assign twiddle4_2_339_imag = T13490 + T13488;
  assign T13488 = $signed(T13489) / $signed(22'h100000);
  assign T13489 = $signed(31'h37e0c9c2) * $signed(16'hffff);
  assign T13490 = {T13493, T13491};
  assign T13491 = $signed(T13492) / $signed(22'h100000);
  assign T13492 = $signed(30'h20cbfa6a) * $signed(16'h0);
  assign T13493 = T13491[6'h2d:6'h2d];
  assign T13494 = T10817[1'h0:1'h0];
  assign T13495 = T10817[1'h1:1'h1];
  assign T13496 = T13521 ? T13511 : T13497;
  assign T13497 = T13510 ? twiddle4_2_341_imag : twiddle4_2_340_imag;
  assign twiddle4_2_340_imag = T13500 + T13498;
  assign T13498 = $signed(T13499) / $signed(22'h100000);
  assign T13499 = $signed(31'h37af8158) * $signed(16'hffff);
  assign T13500 = {T13503, T13501};
  assign T13501 = $signed(T13502) / $signed(22'h100000);
  assign T13502 = $signed(30'h20745b25) * $signed(16'h0);
  assign T13503 = T13501[6'h2d:6'h2d];
  assign twiddle4_2_341_imag = T13506 + T13504;
  assign T13504 = $signed(T13505) / $signed(22'h100000);
  assign T13505 = $signed(31'h377daf89) * $signed(16'hffff);
  assign T13506 = {T13509, T13507};
  assign T13507 = $signed(T13508) / $signed(22'h100000);
  assign T13508 = $signed(30'h201d09b5) * $signed(16'h0);
  assign T13509 = T13507[6'h2d:6'h2d];
  assign T13510 = T10817[1'h0:1'h0];
  assign T13511 = T13520 ? twiddle4_2_343_imag : twiddle4_2_342_imag;
  assign twiddle4_2_342_imag = T13514 + T13512;
  assign T13512 = $signed(T13513) / $signed(22'h100000);
  assign T13513 = $signed(31'h374b54ce) * $signed(16'hffff);
  assign T13514 = $signed(T13515) / $signed(22'h100000);
  assign T13515 = $signed(31'h5fc606f2) * $signed(16'h0);
  assign twiddle4_2_343_imag = T13518 + T13516;
  assign T13516 = $signed(T13517) / $signed(22'h100000);
  assign T13517 = $signed(31'h371871a4) * $signed(16'hffff);
  assign T13518 = $signed(T13519) / $signed(22'h100000);
  assign T13519 = $signed(31'h5f6f53b3) * $signed(16'h0);
  assign T13520 = T10817[1'h0:1'h0];
  assign T13521 = T10817[1'h1:1'h1];
  assign T13522 = T10817[2'h2:2'h2];
  assign T13523 = T13568 ? T13546 : T13524;
  assign T13524 = T13545 ? T13535 : T13525;
  assign T13525 = T13534 ? twiddle4_2_345_imag : twiddle4_2_344_imag;
  assign twiddle4_2_344_imag = T13528 + T13526;
  assign T13526 = $signed(T13527) / $signed(22'h100000);
  assign T13527 = $signed(31'h36e5068a) * $signed(16'hffff);
  assign T13528 = $signed(T13529) / $signed(22'h100000);
  assign T13529 = $signed(31'h5f18f0ce) * $signed(16'h0);
  assign twiddle4_2_345_imag = T13532 + T13530;
  assign T13530 = $signed(T13531) / $signed(22'h100000);
  assign T13531 = $signed(31'h36b113fd) * $signed(16'hffff);
  assign T13532 = $signed(T13533) / $signed(22'h100000);
  assign T13533 = $signed(31'h5ec2df18) * $signed(16'h0);
  assign T13534 = T10817[1'h0:1'h0];
  assign T13535 = T13544 ? twiddle4_2_347_imag : twiddle4_2_346_imag;
  assign twiddle4_2_346_imag = T13538 + T13536;
  assign T13536 = $signed(T13537) / $signed(22'h100000);
  assign T13537 = $signed(31'h367c9a7d) * $signed(16'hffff);
  assign T13538 = $signed(T13539) / $signed(22'h100000);
  assign T13539 = $signed(31'h5e6d1f66) * $signed(16'h0);
  assign twiddle4_2_347_imag = T13542 + T13540;
  assign T13540 = $signed(T13541) / $signed(22'h100000);
  assign T13541 = $signed(31'h36479a8e) * $signed(16'hffff);
  assign T13542 = $signed(T13543) / $signed(22'h100000);
  assign T13543 = $signed(31'h5e17b28a) * $signed(16'h0);
  assign T13544 = T10817[1'h0:1'h0];
  assign T13545 = T10817[1'h1:1'h1];
  assign T13546 = T13567 ? T13557 : T13547;
  assign T13547 = T13556 ? twiddle4_2_349_imag : twiddle4_2_348_imag;
  assign twiddle4_2_348_imag = T13550 + T13548;
  assign T13548 = $signed(T13549) / $signed(22'h100000);
  assign T13549 = $signed(31'h361214b0) * $signed(16'hffff);
  assign T13550 = $signed(T13551) / $signed(22'h100000);
  assign T13551 = $signed(31'h5dc29958) * $signed(16'h0);
  assign twiddle4_2_349_imag = T13554 + T13552;
  assign T13552 = $signed(T13553) / $signed(22'h100000);
  assign T13553 = $signed(31'h35dc0968) * $signed(16'hffff);
  assign T13554 = $signed(T13555) / $signed(22'h100000);
  assign T13555 = $signed(31'h5d6dd4a2) * $signed(16'h0);
  assign T13556 = T10817[1'h0:1'h0];
  assign T13557 = T13566 ? twiddle4_2_351_imag : twiddle4_2_350_imag;
  assign twiddle4_2_350_imag = T13560 + T13558;
  assign T13558 = $signed(T13559) / $signed(22'h100000);
  assign T13559 = $signed(31'h35a5793c) * $signed(16'hffff);
  assign T13560 = $signed(T13561) / $signed(22'h100000);
  assign T13561 = $signed(31'h5d196539) * $signed(16'h0);
  assign twiddle4_2_351_imag = T13564 + T13562;
  assign T13562 = $signed(T13563) / $signed(22'h100000);
  assign T13563 = $signed(31'h356e64b2) * $signed(16'hffff);
  assign T13564 = $signed(T13565) / $signed(22'h100000);
  assign T13565 = $signed(31'h5cc54bed) * $signed(16'h0);
  assign T13566 = T10817[1'h0:1'h0];
  assign T13567 = T10817[1'h1:1'h1];
  assign T13568 = T10817[2'h2:2'h2];
  assign T13569 = T10817[2'h3:2'h3];
  assign T13570 = T10817[3'h4:3'h4];
  assign T13571 = T13760 ? T13666 : T13572;
  assign T13572 = T13665 ? T13619 : T13573;
  assign T13573 = T13618 ? T13596 : T13574;
  assign T13574 = T13595 ? T13585 : T13575;
  assign T13575 = T13584 ? twiddle4_2_353_imag : twiddle4_2_352_imag;
  assign twiddle4_2_352_imag = T13578 + T13576;
  assign T13576 = $signed(T13577) / $signed(22'h100000);
  assign T13577 = $signed(31'h3536cc52) * $signed(16'hffff);
  assign T13578 = $signed(T13579) / $signed(22'h100000);
  assign T13579 = $signed(31'h5c71898d) * $signed(16'h0);
  assign twiddle4_2_353_imag = T13582 + T13580;
  assign T13580 = $signed(T13581) / $signed(22'h100000);
  assign T13581 = $signed(31'h34feb0a5) * $signed(16'hffff);
  assign T13582 = $signed(T13583) / $signed(22'h100000);
  assign T13583 = $signed(31'h5c1e1ee9) * $signed(16'h0);
  assign T13584 = T10817[1'h0:1'h0];
  assign T13585 = T13594 ? twiddle4_2_355_imag : twiddle4_2_354_imag;
  assign twiddle4_2_354_imag = T13588 + T13586;
  assign T13586 = $signed(T13587) / $signed(22'h100000);
  assign T13587 = $signed(31'h34c61236) * $signed(16'hffff);
  assign T13588 = $signed(T13589) / $signed(22'h100000);
  assign T13589 = $signed(31'h5bcb0cce) * $signed(16'h0);
  assign twiddle4_2_355_imag = T13592 + T13590;
  assign T13590 = $signed(T13591) / $signed(22'h100000);
  assign T13591 = $signed(31'h348cf190) * $signed(16'hffff);
  assign T13592 = $signed(T13593) / $signed(22'h100000);
  assign T13593 = $signed(31'h5b785409) * $signed(16'h0);
  assign T13594 = T10817[1'h0:1'h0];
  assign T13595 = T10817[1'h1:1'h1];
  assign T13596 = T13617 ? T13607 : T13597;
  assign T13597 = T13606 ? twiddle4_2_357_imag : twiddle4_2_356_imag;
  assign twiddle4_2_356_imag = T13600 + T13598;
  assign T13598 = $signed(T13599) / $signed(22'h100000);
  assign T13599 = $signed(31'h34534f40) * $signed(16'hffff);
  assign T13600 = $signed(T13601) / $signed(22'h100000);
  assign T13601 = $signed(31'h5b25f567) * $signed(16'h0);
  assign twiddle4_2_357_imag = T13604 + T13602;
  assign T13602 = $signed(T13603) / $signed(22'h100000);
  assign T13603 = $signed(31'h34192bd5) * $signed(16'hffff);
  assign T13604 = $signed(T13605) / $signed(22'h100000);
  assign T13605 = $signed(31'h5ad3f1b2) * $signed(16'h0);
  assign T13606 = T10817[1'h0:1'h0];
  assign T13607 = T13616 ? twiddle4_2_359_imag : twiddle4_2_358_imag;
  assign twiddle4_2_358_imag = T13610 + T13608;
  assign T13608 = $signed(T13609) / $signed(22'h100000);
  assign T13609 = $signed(31'h33de87de) * $signed(16'hffff);
  assign T13610 = $signed(T13611) / $signed(22'h100000);
  assign T13611 = $signed(31'h5a8249b5) * $signed(16'h0);
  assign twiddle4_2_359_imag = T13614 + T13612;
  assign T13612 = $signed(T13613) / $signed(22'h100000);
  assign T13613 = $signed(31'h33a363eb) * $signed(16'hffff);
  assign T13614 = $signed(T13615) / $signed(22'h100000);
  assign T13615 = $signed(31'h5a30fe39) * $signed(16'h0);
  assign T13616 = T10817[1'h0:1'h0];
  assign T13617 = T10817[1'h1:1'h1];
  assign T13618 = T10817[2'h2:2'h2];
  assign T13619 = T13664 ? T13642 : T13620;
  assign T13620 = T13641 ? T13631 : T13621;
  assign T13621 = T13630 ? twiddle4_2_361_imag : twiddle4_2_360_imag;
  assign twiddle4_2_360_imag = T13624 + T13622;
  assign T13622 = $signed(T13623) / $signed(22'h100000);
  assign T13623 = $signed(31'h3367c08f) * $signed(16'hffff);
  assign T13624 = $signed(T13625) / $signed(22'h100000);
  assign T13625 = $signed(31'h59e01007) * $signed(16'h0);
  assign twiddle4_2_361_imag = T13628 + T13626;
  assign T13626 = $signed(T13627) / $signed(22'h100000);
  assign T13627 = $signed(31'h332b9e5d) * $signed(16'hffff);
  assign T13628 = $signed(T13629) / $signed(22'h100000);
  assign T13629 = $signed(31'h598f7fe6) * $signed(16'h0);
  assign T13630 = T10817[1'h0:1'h0];
  assign T13631 = T13640 ? twiddle4_2_363_imag : twiddle4_2_362_imag;
  assign twiddle4_2_362_imag = T13634 + T13632;
  assign T13632 = $signed(T13633) / $signed(22'h100000);
  assign T13633 = $signed(31'h32eefde9) * $signed(16'hffff);
  assign T13634 = $signed(T13635) / $signed(22'h100000);
  assign T13635 = $signed(31'h593f4e9e) * $signed(16'h0);
  assign twiddle4_2_363_imag = T13638 + T13636;
  assign T13636 = $signed(T13637) / $signed(22'h100000);
  assign T13637 = $signed(31'h32b1dfc9) * $signed(16'hffff);
  assign T13638 = $signed(T13639) / $signed(22'h100000);
  assign T13639 = $signed(31'h58ef7cf5) * $signed(16'h0);
  assign T13640 = T10817[1'h0:1'h0];
  assign T13641 = T10817[1'h1:1'h1];
  assign T13642 = T13663 ? T13653 : T13643;
  assign T13643 = T13652 ? twiddle4_2_365_imag : twiddle4_2_364_imag;
  assign twiddle4_2_364_imag = T13646 + T13644;
  assign T13644 = $signed(T13645) / $signed(22'h100000);
  assign T13645 = $signed(31'h32744493) * $signed(16'hffff);
  assign T13646 = $signed(T13647) / $signed(22'h100000);
  assign T13647 = $signed(31'h58a00bae) * $signed(16'h0);
  assign twiddle4_2_365_imag = T13650 + T13648;
  assign T13648 = $signed(T13649) / $signed(22'h100000);
  assign T13649 = $signed(31'h32362cdf) * $signed(16'hffff);
  assign T13650 = $signed(T13651) / $signed(22'h100000);
  assign T13651 = $signed(31'h5850fb8f) * $signed(16'h0);
  assign T13652 = T10817[1'h0:1'h0];
  assign T13653 = T13662 ? twiddle4_2_367_imag : twiddle4_2_366_imag;
  assign twiddle4_2_366_imag = T13656 + T13654;
  assign T13654 = $signed(T13655) / $signed(22'h100000);
  assign T13655 = $signed(31'h31f79947) * $signed(16'hffff);
  assign T13656 = $signed(T13657) / $signed(22'h100000);
  assign T13657 = $signed(31'h58024d5a) * $signed(16'h0);
  assign twiddle4_2_367_imag = T13660 + T13658;
  assign T13658 = $signed(T13659) / $signed(22'h100000);
  assign T13659 = $signed(31'h31b88a66) * $signed(16'hffff);
  assign T13660 = $signed(T13661) / $signed(22'h100000);
  assign T13661 = $signed(31'h57b401d1) * $signed(16'h0);
  assign T13662 = T10817[1'h0:1'h0];
  assign T13663 = T10817[1'h1:1'h1];
  assign T13664 = T10817[2'h2:2'h2];
  assign T13665 = T10817[2'h3:2'h3];
  assign T13666 = T13759 ? T13713 : T13667;
  assign T13667 = T13712 ? T13690 : T13668;
  assign T13668 = T13689 ? T13679 : T13669;
  assign T13669 = T13678 ? twiddle4_2_369_imag : twiddle4_2_368_imag;
  assign twiddle4_2_368_imag = T13672 + T13670;
  assign T13670 = $signed(T13671) / $signed(22'h100000);
  assign T13671 = $signed(31'h317900d6) * $signed(16'hffff);
  assign T13672 = $signed(T13673) / $signed(22'h100000);
  assign T13673 = $signed(31'h576619b6) * $signed(16'h0);
  assign twiddle4_2_369_imag = T13676 + T13674;
  assign T13674 = $signed(T13675) / $signed(22'h100000);
  assign T13675 = $signed(31'h3138fd34) * $signed(16'hffff);
  assign T13676 = $signed(T13677) / $signed(22'h100000);
  assign T13677 = $signed(31'h571895c9) * $signed(16'h0);
  assign T13678 = T10817[1'h0:1'h0];
  assign T13679 = T13688 ? twiddle4_2_371_imag : twiddle4_2_370_imag;
  assign twiddle4_2_370_imag = T13682 + T13680;
  assign T13680 = $signed(T13681) / $signed(22'h100000);
  assign T13681 = $signed(31'h30f8801f) * $signed(16'hffff);
  assign T13682 = $signed(T13683) / $signed(22'h100000);
  assign T13683 = $signed(31'h56cb76c9) * $signed(16'h0);
  assign twiddle4_2_371_imag = T13686 + T13684;
  assign T13684 = $signed(T13685) / $signed(22'h100000);
  assign T13685 = $signed(31'h30b78a35) * $signed(16'hffff);
  assign T13686 = $signed(T13687) / $signed(22'h100000);
  assign T13687 = $signed(31'h567ebd75) * $signed(16'h0);
  assign T13688 = T10817[1'h0:1'h0];
  assign T13689 = T10817[1'h1:1'h1];
  assign T13690 = T13711 ? T13701 : T13691;
  assign T13691 = T13700 ? twiddle4_2_373_imag : twiddle4_2_372_imag;
  assign twiddle4_2_372_imag = T13694 + T13692;
  assign T13692 = $signed(T13693) / $signed(22'h100000);
  assign T13693 = $signed(31'h30761c17) * $signed(16'hffff);
  assign T13694 = $signed(T13695) / $signed(22'h100000);
  assign T13695 = $signed(31'h56326a89) * $signed(16'h0);
  assign twiddle4_2_373_imag = T13698 + T13696;
  assign T13696 = $signed(T13697) / $signed(22'h100000);
  assign T13697 = $signed(31'h30343667) * $signed(16'hffff);
  assign T13698 = $signed(T13699) / $signed(22'h100000);
  assign T13699 = $signed(31'h55e67ec2) * $signed(16'h0);
  assign T13700 = T10817[1'h0:1'h0];
  assign T13701 = T13710 ? twiddle4_2_375_imag : twiddle4_2_374_imag;
  assign twiddle4_2_374_imag = T13704 + T13702;
  assign T13702 = $signed(T13703) / $signed(22'h100000);
  assign T13703 = $signed(31'h2ff1d9c6) * $signed(16'hffff);
  assign T13704 = $signed(T13705) / $signed(22'h100000);
  assign T13705 = $signed(31'h559afadb) * $signed(16'h0);
  assign twiddle4_2_375_imag = T13708 + T13706;
  assign T13706 = $signed(T13707) / $signed(22'h100000);
  assign T13707 = $signed(31'h2faf06d9) * $signed(16'hffff);
  assign T13708 = $signed(T13709) / $signed(22'h100000);
  assign T13709 = $signed(31'h554fdf8f) * $signed(16'h0);
  assign T13710 = T10817[1'h0:1'h0];
  assign T13711 = T10817[1'h1:1'h1];
  assign T13712 = T10817[2'h2:2'h2];
  assign T13713 = T13758 ? T13736 : T13714;
  assign T13714 = T13735 ? T13725 : T13715;
  assign T13715 = T13724 ? twiddle4_2_377_imag : twiddle4_2_376_imag;
  assign twiddle4_2_376_imag = T13718 + T13716;
  assign T13716 = $signed(T13717) / $signed(22'h100000);
  assign T13717 = $signed(31'h2f6bbe44) * $signed(16'hffff);
  assign T13718 = $signed(T13719) / $signed(22'h100000);
  assign T13719 = $signed(31'h55052d97) * $signed(16'h0);
  assign twiddle4_2_377_imag = T13722 + T13720;
  assign T13720 = $signed(T13721) / $signed(22'h100000);
  assign T13721 = $signed(31'h2f2800ae) * $signed(16'hffff);
  assign T13722 = $signed(T13723) / $signed(22'h100000);
  assign T13723 = $signed(31'h54bae5ac) * $signed(16'h0);
  assign T13724 = T10817[1'h0:1'h0];
  assign T13725 = T13734 ? twiddle4_2_379_imag : twiddle4_2_378_imag;
  assign twiddle4_2_378_imag = T13728 + T13726;
  assign T13726 = $signed(T13727) / $signed(22'h100000);
  assign T13727 = $signed(31'h2ee3cebe) * $signed(16'hffff);
  assign T13728 = $signed(T13729) / $signed(22'h100000);
  assign T13729 = $signed(31'h54710884) * $signed(16'h0);
  assign twiddle4_2_379_imag = T13732 + T13730;
  assign T13730 = $signed(T13731) / $signed(22'h100000);
  assign T13731 = $signed(31'h2e9f291b) * $signed(16'hffff);
  assign T13732 = $signed(T13733) / $signed(22'h100000);
  assign T13733 = $signed(31'h542796d5) * $signed(16'h0);
  assign T13734 = T10817[1'h0:1'h0];
  assign T13735 = T10817[1'h1:1'h1];
  assign T13736 = T13757 ? T13747 : T13737;
  assign T13737 = T13746 ? twiddle4_2_381_imag : twiddle4_2_380_imag;
  assign twiddle4_2_380_imag = T13740 + T13738;
  assign T13738 = $signed(T13739) / $signed(22'h100000);
  assign T13739 = $signed(31'h2e5a106f) * $signed(16'hffff);
  assign T13740 = $signed(T13741) / $signed(22'h100000);
  assign T13741 = $signed(31'h53de9156) * $signed(16'h0);
  assign twiddle4_2_381_imag = T13744 + T13742;
  assign T13742 = $signed(T13743) / $signed(22'h100000);
  assign T13743 = $signed(31'h2e148566) * $signed(16'hffff);
  assign T13744 = $signed(T13745) / $signed(22'h100000);
  assign T13745 = $signed(31'h5395f8ba) * $signed(16'h0);
  assign T13746 = T10817[1'h0:1'h0];
  assign T13747 = T13756 ? twiddle4_2_383_imag : twiddle4_2_382_imag;
  assign twiddle4_2_382_imag = T13750 + T13748;
  assign T13748 = $signed(T13749) / $signed(22'h100000);
  assign T13749 = $signed(31'h2dce88a9) * $signed(16'hffff);
  assign T13750 = $signed(T13751) / $signed(22'h100000);
  assign T13751 = $signed(31'h534dcdb5) * $signed(16'h0);
  assign twiddle4_2_383_imag = T13754 + T13752;
  assign T13752 = $signed(T13753) / $signed(22'h100000);
  assign T13753 = $signed(31'h2d881ae7) * $signed(16'hffff);
  assign T13754 = $signed(T13755) / $signed(22'h100000);
  assign T13755 = $signed(31'h530610f7) * $signed(16'h0);
  assign T13756 = T10817[1'h0:1'h0];
  assign T13757 = T10817[1'h1:1'h1];
  assign T13758 = T10817[2'h2:2'h2];
  assign T13759 = T10817[2'h3:2'h3];
  assign T13760 = T10817[3'h4:3'h4];
  assign T13761 = T10817[3'h5:3'h5];
  assign T13762 = T13336[6'h2e:6'h2e];
  assign T13763 = T10817[3'h6:3'h6];
  assign T13764 = {T14742, T13765};
  assign T13765 = T14741 ? T14190 : T13766;
  assign T13766 = T14189 ? T13957 : T13767;
  assign T13767 = T13956 ? T13862 : T13768;
  assign T13768 = T13861 ? T13815 : T13769;
  assign T13769 = T13814 ? T13792 : T13770;
  assign T13770 = T13791 ? T13781 : T13771;
  assign T13771 = T13780 ? twiddle4_2_385_imag : twiddle4_2_384_imag;
  assign twiddle4_2_384_imag = T13774 + T13772;
  assign T13772 = $signed(T13773) / $signed(22'h100000);
  assign T13773 = $signed(31'h2d413ccc) * $signed(16'hffff);
  assign T13774 = $signed(T13775) / $signed(22'h100000);
  assign T13775 = $signed(31'h52bec334) * $signed(16'h0);
  assign twiddle4_2_385_imag = T13778 + T13776;
  assign T13776 = $signed(T13777) / $signed(22'h100000);
  assign T13777 = $signed(31'h2cf9ef09) * $signed(16'hffff);
  assign T13778 = $signed(T13779) / $signed(22'h100000);
  assign T13779 = $signed(31'h5277e519) * $signed(16'h0);
  assign T13780 = T10817[1'h0:1'h0];
  assign T13781 = T13790 ? twiddle4_2_387_imag : twiddle4_2_386_imag;
  assign twiddle4_2_386_imag = T13784 + T13782;
  assign T13782 = $signed(T13783) / $signed(22'h100000);
  assign T13783 = $signed(31'h2cb2324b) * $signed(16'hffff);
  assign T13784 = $signed(T13785) / $signed(22'h100000);
  assign T13785 = $signed(31'h52317757) * $signed(16'h0);
  assign twiddle4_2_387_imag = T13788 + T13786;
  assign T13786 = $signed(T13787) / $signed(22'h100000);
  assign T13787 = $signed(31'h2c6a0746) * $signed(16'hffff);
  assign T13788 = $signed(T13789) / $signed(22'h100000);
  assign T13789 = $signed(31'h51eb7a9a) * $signed(16'h0);
  assign T13790 = T10817[1'h0:1'h0];
  assign T13791 = T10817[1'h1:1'h1];
  assign T13792 = T13813 ? T13803 : T13793;
  assign T13793 = T13802 ? twiddle4_2_389_imag : twiddle4_2_388_imag;
  assign twiddle4_2_388_imag = T13796 + T13794;
  assign T13794 = $signed(T13795) / $signed(22'h100000);
  assign T13795 = $signed(31'h2c216eaa) * $signed(16'hffff);
  assign T13796 = $signed(T13797) / $signed(22'h100000);
  assign T13797 = $signed(31'h51a5ef91) * $signed(16'h0);
  assign twiddle4_2_389_imag = T13800 + T13798;
  assign T13798 = $signed(T13799) / $signed(22'h100000);
  assign T13799 = $signed(31'h2bd8692b) * $signed(16'hffff);
  assign T13800 = $signed(T13801) / $signed(22'h100000);
  assign T13801 = $signed(31'h5160d6e5) * $signed(16'h0);
  assign T13802 = T10817[1'h0:1'h0];
  assign T13803 = T13812 ? twiddle4_2_391_imag : twiddle4_2_390_imag;
  assign twiddle4_2_390_imag = T13806 + T13804;
  assign T13804 = $signed(T13805) / $signed(22'h100000);
  assign T13805 = $signed(31'h2b8ef77c) * $signed(16'hffff);
  assign T13806 = $signed(T13807) / $signed(22'h100000);
  assign T13807 = $signed(31'h511c3142) * $signed(16'h0);
  assign twiddle4_2_391_imag = T13810 + T13808;
  assign T13808 = $signed(T13809) / $signed(22'h100000);
  assign T13809 = $signed(31'h2b451a54) * $signed(16'hffff);
  assign T13810 = $signed(T13811) / $signed(22'h100000);
  assign T13811 = $signed(31'h50d7ff52) * $signed(16'h0);
  assign T13812 = T10817[1'h0:1'h0];
  assign T13813 = T10817[1'h1:1'h1];
  assign T13814 = T10817[2'h2:2'h2];
  assign T13815 = T13860 ? T13838 : T13816;
  assign T13816 = T13837 ? T13827 : T13817;
  assign T13817 = T13826 ? twiddle4_2_393_imag : twiddle4_2_392_imag;
  assign twiddle4_2_392_imag = T13820 + T13818;
  assign T13818 = $signed(T13819) / $signed(22'h100000);
  assign T13819 = $signed(31'h2afad269) * $signed(16'hffff);
  assign T13820 = $signed(T13821) / $signed(22'h100000);
  assign T13821 = $signed(31'h509441bc) * $signed(16'h0);
  assign twiddle4_2_393_imag = T13824 + T13822;
  assign T13822 = $signed(T13823) / $signed(22'h100000);
  assign T13823 = $signed(31'h2ab02071) * $signed(16'hffff);
  assign T13824 = $signed(T13825) / $signed(22'h100000);
  assign T13825 = $signed(31'h5050f927) * $signed(16'h0);
  assign T13826 = T10817[1'h0:1'h0];
  assign T13827 = T13836 ? twiddle4_2_395_imag : twiddle4_2_394_imag;
  assign twiddle4_2_394_imag = T13830 + T13828;
  assign T13828 = $signed(T13829) / $signed(22'h100000);
  assign T13829 = $signed(31'h2a650525) * $signed(16'hffff);
  assign T13830 = $signed(T13831) / $signed(22'h100000);
  assign T13831 = $signed(31'h500e263a) * $signed(16'h0);
  assign twiddle4_2_395_imag = T13834 + T13832;
  assign T13832 = $signed(T13833) / $signed(22'h100000);
  assign T13833 = $signed(31'h2a19813e) * $signed(16'hffff);
  assign T13834 = $signed(T13835) / $signed(22'h100000);
  assign T13835 = $signed(31'h4fcbc999) * $signed(16'h0);
  assign T13836 = T10817[1'h0:1'h0];
  assign T13837 = T10817[1'h1:1'h1];
  assign T13838 = T13859 ? T13849 : T13839;
  assign T13839 = T13848 ? twiddle4_2_397_imag : twiddle4_2_396_imag;
  assign twiddle4_2_396_imag = T13842 + T13840;
  assign T13840 = $signed(T13841) / $signed(22'h100000);
  assign T13841 = $signed(31'h29cd9577) * $signed(16'hffff);
  assign T13842 = $signed(T13843) / $signed(22'h100000);
  assign T13843 = $signed(31'h4f89e3e9) * $signed(16'h0);
  assign twiddle4_2_397_imag = T13846 + T13844;
  assign T13844 = $signed(T13845) / $signed(22'h100000);
  assign T13845 = $signed(31'h2981428b) * $signed(16'hffff);
  assign T13846 = $signed(T13847) / $signed(22'h100000);
  assign T13847 = $signed(31'h4f4875cb) * $signed(16'h0);
  assign T13848 = T10817[1'h0:1'h0];
  assign T13849 = T13858 ? twiddle4_2_399_imag : twiddle4_2_398_imag;
  assign twiddle4_2_398_imag = T13852 + T13850;
  assign T13850 = $signed(T13851) / $signed(22'h100000);
  assign T13851 = $signed(31'h29348937) * $signed(16'hffff);
  assign T13852 = $signed(T13853) / $signed(22'h100000);
  assign T13853 = $signed(31'h4f077fe1) * $signed(16'h0);
  assign twiddle4_2_399_imag = T13856 + T13854;
  assign T13854 = $signed(T13855) / $signed(22'h100000);
  assign T13855 = $signed(31'h28e76a37) * $signed(16'hffff);
  assign T13856 = $signed(T13857) / $signed(22'h100000);
  assign T13857 = $signed(31'h4ec702cc) * $signed(16'h0);
  assign T13858 = T10817[1'h0:1'h0];
  assign T13859 = T10817[1'h1:1'h1];
  assign T13860 = T10817[2'h2:2'h2];
  assign T13861 = T10817[2'h3:2'h3];
  assign T13862 = T13955 ? T13909 : T13863;
  assign T13863 = T13908 ? T13886 : T13864;
  assign T13864 = T13885 ? T13875 : T13865;
  assign T13865 = T13874 ? twiddle4_2_401_imag : twiddle4_2_400_imag;
  assign twiddle4_2_400_imag = T13868 + T13866;
  assign T13866 = $signed(T13867) / $signed(22'h100000);
  assign T13867 = $signed(31'h2899e64a) * $signed(16'hffff);
  assign T13868 = $signed(T13869) / $signed(22'h100000);
  assign T13869 = $signed(31'h4e86ff2a) * $signed(16'h0);
  assign twiddle4_2_401_imag = T13872 + T13870;
  assign T13870 = $signed(T13871) / $signed(22'h100000);
  assign T13871 = $signed(31'h284bfe2f) * $signed(16'hffff);
  assign T13872 = $signed(T13873) / $signed(22'h100000);
  assign T13873 = $signed(31'h4e47759a) * $signed(16'h0);
  assign T13874 = T10817[1'h0:1'h0];
  assign T13875 = T13884 ? twiddle4_2_403_imag : twiddle4_2_402_imag;
  assign twiddle4_2_402_imag = T13878 + T13876;
  assign T13876 = $signed(T13877) / $signed(22'h100000);
  assign T13877 = $signed(31'h27fdb2a6) * $signed(16'hffff);
  assign T13878 = $signed(T13879) / $signed(22'h100000);
  assign T13879 = $signed(31'h4e0866b9) * $signed(16'h0);
  assign twiddle4_2_403_imag = T13882 + T13880;
  assign T13880 = $signed(T13881) / $signed(22'h100000);
  assign T13881 = $signed(31'h27af0471) * $signed(16'hffff);
  assign T13882 = $signed(T13883) / $signed(22'h100000);
  assign T13883 = $signed(31'h4dc9d321) * $signed(16'h0);
  assign T13884 = T10817[1'h0:1'h0];
  assign T13885 = T10817[1'h1:1'h1];
  assign T13886 = T13907 ? T13897 : T13887;
  assign T13887 = T13896 ? twiddle4_2_405_imag : twiddle4_2_404_imag;
  assign twiddle4_2_404_imag = T13890 + T13888;
  assign T13888 = $signed(T13889) / $signed(22'h100000);
  assign T13889 = $signed(31'h275ff452) * $signed(16'hffff);
  assign T13890 = $signed(T13891) / $signed(22'h100000);
  assign T13891 = $signed(31'h4d8bbb6d) * $signed(16'h0);
  assign twiddle4_2_405_imag = T13894 + T13892;
  assign T13892 = $signed(T13893) / $signed(22'h100000);
  assign T13893 = $signed(31'h2710830b) * $signed(16'hffff);
  assign T13894 = $signed(T13895) / $signed(22'h100000);
  assign T13895 = $signed(31'h4d4e2037) * $signed(16'h0);
  assign T13896 = T10817[1'h0:1'h0];
  assign T13897 = T13906 ? twiddle4_2_407_imag : twiddle4_2_406_imag;
  assign twiddle4_2_406_imag = T13900 + T13898;
  assign T13898 = $signed(T13899) / $signed(22'h100000);
  assign T13899 = $signed(31'h26c0b162) * $signed(16'hffff);
  assign T13900 = $signed(T13901) / $signed(22'h100000);
  assign T13901 = $signed(31'h4d110217) * $signed(16'h0);
  assign twiddle4_2_407_imag = T13904 + T13902;
  assign T13902 = $signed(T13903) / $signed(22'h100000);
  assign T13903 = $signed(31'h2670801a) * $signed(16'hffff);
  assign T13904 = $signed(T13905) / $signed(22'h100000);
  assign T13905 = $signed(31'h4cd461a3) * $signed(16'h0);
  assign T13906 = T10817[1'h0:1'h0];
  assign T13907 = T10817[1'h1:1'h1];
  assign T13908 = T10817[2'h2:2'h2];
  assign T13909 = T13954 ? T13932 : T13910;
  assign T13910 = T13931 ? T13921 : T13911;
  assign T13911 = T13920 ? twiddle4_2_409_imag : twiddle4_2_408_imag;
  assign twiddle4_2_408_imag = T13914 + T13912;
  assign T13912 = $signed(T13913) / $signed(22'h100000);
  assign T13913 = $signed(31'h261feff9) * $signed(16'hffff);
  assign T13914 = $signed(T13915) / $signed(22'h100000);
  assign T13915 = $signed(31'h4c983f71) * $signed(16'h0);
  assign twiddle4_2_409_imag = T13918 + T13916;
  assign T13916 = $signed(T13917) / $signed(22'h100000);
  assign T13917 = $signed(31'h25cf01c7) * $signed(16'hffff);
  assign T13918 = $signed(T13919) / $signed(22'h100000);
  assign T13919 = $signed(31'h4c5c9c15) * $signed(16'h0);
  assign T13920 = T10817[1'h0:1'h0];
  assign T13921 = T13930 ? twiddle4_2_411_imag : twiddle4_2_410_imag;
  assign twiddle4_2_410_imag = T13924 + T13922;
  assign T13922 = $signed(T13923) / $signed(22'h100000);
  assign T13923 = $signed(31'h257db64b) * $signed(16'hffff);
  assign T13924 = $signed(T13925) / $signed(22'h100000);
  assign T13925 = $signed(31'h4c217822) * $signed(16'h0);
  assign twiddle4_2_411_imag = T13928 + T13926;
  assign T13926 = $signed(T13927) / $signed(22'h100000);
  assign T13927 = $signed(31'h252c0e4e) * $signed(16'hffff);
  assign T13928 = $signed(T13929) / $signed(22'h100000);
  assign T13929 = $signed(31'h4be6d42b) * $signed(16'h0);
  assign T13930 = T10817[1'h0:1'h0];
  assign T13931 = T10817[1'h1:1'h1];
  assign T13932 = T13953 ? T13943 : T13933;
  assign T13933 = T13942 ? twiddle4_2_413_imag : twiddle4_2_412_imag;
  assign twiddle4_2_412_imag = T13936 + T13934;
  assign T13934 = $signed(T13935) / $signed(22'h100000);
  assign T13935 = $signed(31'h24da0a99) * $signed(16'hffff);
  assign T13936 = $signed(T13937) / $signed(22'h100000);
  assign T13937 = $signed(31'h4bacb0c0) * $signed(16'h0);
  assign twiddle4_2_413_imag = T13940 + T13938;
  assign T13938 = $signed(T13939) / $signed(22'h100000);
  assign T13939 = $signed(31'h2487abf7) * $signed(16'hffff);
  assign T13940 = $signed(T13941) / $signed(22'h100000);
  assign T13941 = $signed(31'h4b730e70) * $signed(16'h0);
  assign T13942 = T10817[1'h0:1'h0];
  assign T13943 = T13952 ? twiddle4_2_415_imag : twiddle4_2_414_imag;
  assign twiddle4_2_414_imag = T13946 + T13944;
  assign T13944 = $signed(T13945) / $signed(22'h100000);
  assign T13945 = $signed(31'h2434f332) * $signed(16'hffff);
  assign T13946 = $signed(T13947) / $signed(22'h100000);
  assign T13947 = $signed(31'h4b39edca) * $signed(16'h0);
  assign twiddle4_2_415_imag = T13950 + T13948;
  assign T13948 = $signed(T13949) / $signed(22'h100000);
  assign T13949 = $signed(31'h23e1e117) * $signed(16'hffff);
  assign T13950 = $signed(T13951) / $signed(22'h100000);
  assign T13951 = $signed(31'h4b014f5b) * $signed(16'h0);
  assign T13952 = T10817[1'h0:1'h0];
  assign T13953 = T10817[1'h1:1'h1];
  assign T13954 = T10817[2'h2:2'h2];
  assign T13955 = T10817[2'h3:2'h3];
  assign T13956 = T10817[3'h4:3'h4];
  assign T13957 = T14188 ? T14062 : T13958;
  assign T13958 = T14061 ? T14005 : T13959;
  assign T13959 = T14004 ? T13982 : T13960;
  assign T13960 = T13981 ? T13971 : T13961;
  assign T13961 = T13970 ? twiddle4_2_417_imag : twiddle4_2_416_imag;
  assign twiddle4_2_416_imag = T13964 + T13962;
  assign T13962 = $signed(T13963) / $signed(22'h100000);
  assign T13963 = $signed(31'h238e7673) * $signed(16'hffff);
  assign T13964 = $signed(T13965) / $signed(22'h100000);
  assign T13965 = $signed(31'h4ac933ae) * $signed(16'h0);
  assign twiddle4_2_417_imag = T13968 + T13966;
  assign T13966 = $signed(T13967) / $signed(22'h100000);
  assign T13967 = $signed(31'h233ab413) * $signed(16'hffff);
  assign T13968 = $signed(T13969) / $signed(22'h100000);
  assign T13969 = $signed(31'h4a919b4e) * $signed(16'h0);
  assign T13970 = T10817[1'h0:1'h0];
  assign T13971 = T13980 ? twiddle4_2_419_imag : twiddle4_2_418_imag;
  assign twiddle4_2_418_imag = T13974 + T13972;
  assign T13972 = $signed(T13973) / $signed(22'h100000);
  assign T13973 = $signed(31'h22e69ac7) * $signed(16'hffff);
  assign T13974 = $signed(T13975) / $signed(22'h100000);
  assign T13975 = $signed(31'h4a5a86c4) * $signed(16'h0);
  assign twiddle4_2_419_imag = T13978 + T13976;
  assign T13976 = $signed(T13977) / $signed(22'h100000);
  assign T13977 = $signed(31'h22922b5e) * $signed(16'hffff);
  assign T13978 = $signed(T13979) / $signed(22'h100000);
  assign T13979 = $signed(31'h4a23f698) * $signed(16'h0);
  assign T13980 = T10817[1'h0:1'h0];
  assign T13981 = T10817[1'h1:1'h1];
  assign T13982 = T14003 ? T13993 : T13983;
  assign T13983 = T13992 ? twiddle4_2_421_imag : twiddle4_2_420_imag;
  assign twiddle4_2_420_imag = T13986 + T13984;
  assign T13984 = $signed(T13985) / $signed(22'h100000);
  assign T13985 = $signed(31'h223d66a8) * $signed(16'hffff);
  assign T13986 = $signed(T13987) / $signed(22'h100000);
  assign T13987 = $signed(31'h49edeb50) * $signed(16'h0);
  assign twiddle4_2_421_imag = T13990 + T13988;
  assign T13988 = $signed(T13989) / $signed(22'h100000);
  assign T13989 = $signed(31'h21e84d76) * $signed(16'hffff);
  assign T13990 = $signed(T13991) / $signed(22'h100000);
  assign T13991 = $signed(31'h49b86572) * $signed(16'h0);
  assign T13992 = T10817[1'h0:1'h0];
  assign T13993 = T14002 ? twiddle4_2_423_imag : twiddle4_2_422_imag;
  assign twiddle4_2_422_imag = T13996 + T13994;
  assign T13994 = $signed(T13995) / $signed(22'h100000);
  assign T13995 = $signed(31'h2192e09a) * $signed(16'hffff);
  assign T13996 = $signed(T13997) / $signed(22'h100000);
  assign T13997 = $signed(31'h49836583) * $signed(16'h0);
  assign twiddle4_2_423_imag = T14000 + T13998;
  assign T13998 = $signed(T13999) / $signed(22'h100000);
  assign T13999 = $signed(31'h213d20e8) * $signed(16'hffff);
  assign T14000 = $signed(T14001) / $signed(22'h100000);
  assign T14001 = $signed(31'h494eec03) * $signed(16'h0);
  assign T14002 = T10817[1'h0:1'h0];
  assign T14003 = T10817[1'h1:1'h1];
  assign T14004 = T10817[2'h2:2'h2];
  assign T14005 = T14060 ? T14030 : T14006;
  assign T14006 = T14029 ? T14017 : T14007;
  assign T14007 = T14016 ? twiddle4_2_425_imag : twiddle4_2_424_imag;
  assign twiddle4_2_424_imag = T14010 + T14008;
  assign T14008 = $signed(T14009) / $signed(22'h100000);
  assign T14009 = $signed(31'h20e70f32) * $signed(16'hffff);
  assign T14010 = $signed(T14011) / $signed(22'h100000);
  assign T14011 = $signed(31'h491af976) * $signed(16'h0);
  assign twiddle4_2_425_imag = T14014 + T14012;
  assign T14012 = $signed(T14013) / $signed(22'h100000);
  assign T14013 = $signed(31'h2090ac4d) * $signed(16'hffff);
  assign T14014 = $signed(T14015) / $signed(22'h100000);
  assign T14015 = $signed(31'h48e78e5c) * $signed(16'h0);
  assign T14016 = T10817[1'h0:1'h0];
  assign T14017 = T14028 ? twiddle4_2_427_imag : twiddle4_2_426_imag;
  assign twiddle4_2_426_imag = T14020 + T14018;
  assign T14018 = $signed(T14019) / $signed(22'h100000);
  assign T14019 = $signed(31'h2039f90e) * $signed(16'hffff);
  assign T14020 = $signed(T14021) / $signed(22'h100000);
  assign T14021 = $signed(31'h48b4ab32) * $signed(16'h0);
  assign twiddle4_2_427_imag = T14026 + T14022;
  assign T14022 = {T14025, T14023};
  assign T14023 = $signed(T14024) / $signed(22'h100000);
  assign T14024 = $signed(30'h1fe2f64b) * $signed(16'hffff);
  assign T14025 = T14023[6'h2d:6'h2d];
  assign T14026 = $signed(T14027) / $signed(22'h100000);
  assign T14027 = $signed(31'h48825077) * $signed(16'h0);
  assign T14028 = T10817[1'h0:1'h0];
  assign T14029 = T10817[1'h1:1'h1];
  assign T14030 = T14059 ? T14045 : T14031;
  assign T14031 = T14044 ? twiddle4_2_429_imag : twiddle4_2_428_imag;
  assign twiddle4_2_428_imag = T14036 + T14032;
  assign T14032 = {T14035, T14033};
  assign T14033 = $signed(T14034) / $signed(22'h100000);
  assign T14034 = $signed(30'h1f8ba4db) * $signed(16'hffff);
  assign T14035 = T14033[6'h2d:6'h2d];
  assign T14036 = $signed(T14037) / $signed(22'h100000);
  assign T14037 = $signed(31'h48507ea8) * $signed(16'h0);
  assign twiddle4_2_429_imag = T14042 + T14038;
  assign T14038 = {T14041, T14039};
  assign T14039 = $signed(T14040) / $signed(22'h100000);
  assign T14040 = $signed(30'h1f340596) * $signed(16'hffff);
  assign T14041 = T14039[6'h2d:6'h2d];
  assign T14042 = $signed(T14043) / $signed(22'h100000);
  assign T14043 = $signed(31'h481f363e) * $signed(16'h0);
  assign T14044 = T10817[1'h0:1'h0];
  assign T14045 = T14058 ? twiddle4_2_431_imag : twiddle4_2_430_imag;
  assign twiddle4_2_430_imag = T14050 + T14046;
  assign T14046 = {T14049, T14047};
  assign T14047 = $signed(T14048) / $signed(22'h100000);
  assign T14048 = $signed(30'h1edc1952) * $signed(16'hffff);
  assign T14049 = T14047[6'h2d:6'h2d];
  assign T14050 = $signed(T14051) / $signed(22'h100000);
  assign T14051 = $signed(31'h47ee77b4) * $signed(16'h0);
  assign twiddle4_2_431_imag = T14056 + T14052;
  assign T14052 = {T14055, T14053};
  assign T14053 = $signed(T14054) / $signed(22'h100000);
  assign T14054 = $signed(30'h1e83e0ea) * $signed(16'hffff);
  assign T14055 = T14053[6'h2d:6'h2d];
  assign T14056 = $signed(T14057) / $signed(22'h100000);
  assign T14057 = $signed(31'h47be4381) * $signed(16'h0);
  assign T14058 = T10817[1'h0:1'h0];
  assign T14059 = T10817[1'h1:1'h1];
  assign T14060 = T10817[2'h2:2'h2];
  assign T14061 = T10817[2'h3:2'h3];
  assign T14062 = T14187 ? T14125 : T14063;
  assign T14063 = T14124 ? T14094 : T14064;
  assign T14064 = T14093 ? T14079 : T14065;
  assign T14065 = T14078 ? twiddle4_2_433_imag : twiddle4_2_432_imag;
  assign twiddle4_2_432_imag = T14070 + T14066;
  assign T14066 = {T14069, T14067};
  assign T14067 = $signed(T14068) / $signed(22'h100000);
  assign T14068 = $signed(30'h1e2b5d38) * $signed(16'hffff);
  assign T14069 = T14067[6'h2d:6'h2d];
  assign T14070 = $signed(T14071) / $signed(22'h100000);
  assign T14071 = $signed(31'h478e9a1d) * $signed(16'h0);
  assign twiddle4_2_433_imag = T14076 + T14072;
  assign T14072 = {T14075, T14073};
  assign T14073 = $signed(T14074) / $signed(22'h100000);
  assign T14074 = $signed(30'h1dd28f14) * $signed(16'hffff);
  assign T14075 = T14073[6'h2d:6'h2d];
  assign T14076 = $signed(T14077) / $signed(22'h100000);
  assign T14077 = $signed(31'h475f7bfe) * $signed(16'h0);
  assign T14078 = T10817[1'h0:1'h0];
  assign T14079 = T14092 ? twiddle4_2_435_imag : twiddle4_2_434_imag;
  assign twiddle4_2_434_imag = T14084 + T14080;
  assign T14080 = {T14083, T14081};
  assign T14081 = $signed(T14082) / $signed(22'h100000);
  assign T14082 = $signed(30'h1d79775b) * $signed(16'hffff);
  assign T14083 = T14081[6'h2d:6'h2d];
  assign T14084 = $signed(T14085) / $signed(22'h100000);
  assign T14085 = $signed(31'h4730e997) * $signed(16'h0);
  assign twiddle4_2_435_imag = T14090 + T14086;
  assign T14086 = {T14089, T14087};
  assign T14087 = $signed(T14088) / $signed(22'h100000);
  assign T14088 = $signed(30'h1d2016e8) * $signed(16'hffff);
  assign T14089 = T14087[6'h2d:6'h2d];
  assign T14090 = $signed(T14091) / $signed(22'h100000);
  assign T14091 = $signed(31'h4702e35c) * $signed(16'h0);
  assign T14092 = T10817[1'h0:1'h0];
  assign T14093 = T10817[1'h1:1'h1];
  assign T14094 = T14123 ? T14109 : T14095;
  assign T14095 = T14108 ? twiddle4_2_437_imag : twiddle4_2_436_imag;
  assign twiddle4_2_436_imag = T14100 + T14096;
  assign T14096 = {T14099, T14097};
  assign T14097 = $signed(T14098) / $signed(22'h100000);
  assign T14098 = $signed(30'h1cc66e99) * $signed(16'hffff);
  assign T14099 = T14097[6'h2d:6'h2d];
  assign T14100 = $signed(T14101) / $signed(22'h100000);
  assign T14101 = $signed(31'h46d569be) * $signed(16'h0);
  assign twiddle4_2_437_imag = T14106 + T14102;
  assign T14102 = {T14105, T14103};
  assign T14103 = $signed(T14104) / $signed(22'h100000);
  assign T14104 = $signed(30'h1c6c7f49) * $signed(16'hffff);
  assign T14105 = T14103[6'h2d:6'h2d];
  assign T14106 = $signed(T14107) / $signed(22'h100000);
  assign T14107 = $signed(31'h46a87d2d) * $signed(16'h0);
  assign T14108 = T10817[1'h0:1'h0];
  assign T14109 = T14122 ? twiddle4_2_439_imag : twiddle4_2_438_imag;
  assign twiddle4_2_438_imag = T14114 + T14110;
  assign T14110 = {T14113, T14111};
  assign T14111 = $signed(T14112) / $signed(22'h100000);
  assign T14112 = $signed(30'h1c1249d8) * $signed(16'hffff);
  assign T14113 = T14111[6'h2d:6'h2d];
  assign T14114 = $signed(T14115) / $signed(22'h100000);
  assign T14115 = $signed(31'h467c1e19) * $signed(16'h0);
  assign twiddle4_2_439_imag = T14120 + T14116;
  assign T14116 = {T14119, T14117};
  assign T14117 = $signed(T14118) / $signed(22'h100000);
  assign T14118 = $signed(30'h1bb7cf23) * $signed(16'hffff);
  assign T14119 = T14117[6'h2d:6'h2d];
  assign T14120 = $signed(T14121) / $signed(22'h100000);
  assign T14121 = $signed(31'h46504ced) * $signed(16'h0);
  assign T14122 = T10817[1'h0:1'h0];
  assign T14123 = T10817[1'h1:1'h1];
  assign T14124 = T10817[2'h2:2'h2];
  assign T14125 = T14186 ? T14156 : T14126;
  assign T14126 = T14155 ? T14141 : T14127;
  assign T14127 = T14140 ? twiddle4_2_441_imag : twiddle4_2_440_imag;
  assign twiddle4_2_440_imag = T14132 + T14128;
  assign T14128 = {T14131, T14129};
  assign T14129 = $signed(T14130) / $signed(22'h100000);
  assign T14130 = $signed(30'h1b5d1009) * $signed(16'hffff);
  assign T14131 = T14129[6'h2d:6'h2d];
  assign T14132 = $signed(T14133) / $signed(22'h100000);
  assign T14133 = $signed(31'h46250a18) * $signed(16'h0);
  assign twiddle4_2_441_imag = T14138 + T14134;
  assign T14134 = {T14137, T14135};
  assign T14135 = $signed(T14136) / $signed(22'h100000);
  assign T14136 = $signed(30'h1b020d6c) * $signed(16'hffff);
  assign T14137 = T14135[6'h2d:6'h2d];
  assign T14138 = $signed(T14139) / $signed(22'h100000);
  assign T14139 = $signed(31'h45fa5603) * $signed(16'h0);
  assign T14140 = T10817[1'h0:1'h0];
  assign T14141 = T14154 ? twiddle4_2_443_imag : twiddle4_2_442_imag;
  assign twiddle4_2_442_imag = T14146 + T14142;
  assign T14142 = {T14145, T14143};
  assign T14143 = $signed(T14144) / $signed(22'h100000);
  assign T14144 = $signed(30'h1aa6c82b) * $signed(16'hffff);
  assign T14145 = T14143[6'h2d:6'h2d];
  assign T14146 = $signed(T14147) / $signed(22'h100000);
  assign T14147 = $signed(31'h45d03118) * $signed(16'h0);
  assign twiddle4_2_443_imag = T14152 + T14148;
  assign T14148 = {T14151, T14149};
  assign T14149 = $signed(T14150) / $signed(22'h100000);
  assign T14150 = $signed(30'h1a4b4127) * $signed(16'hffff);
  assign T14151 = T14149[6'h2d:6'h2d];
  assign T14152 = $signed(T14153) / $signed(22'h100000);
  assign T14153 = $signed(31'h45a69bbf) * $signed(16'h0);
  assign T14154 = T10817[1'h0:1'h0];
  assign T14155 = T10817[1'h1:1'h1];
  assign T14156 = T14185 ? T14171 : T14157;
  assign T14157 = T14170 ? twiddle4_2_445_imag : twiddle4_2_444_imag;
  assign twiddle4_2_444_imag = T14162 + T14158;
  assign T14158 = {T14161, T14159};
  assign T14159 = $signed(T14160) / $signed(22'h100000);
  assign T14160 = $signed(30'h19ef7943) * $signed(16'hffff);
  assign T14161 = T14159[6'h2d:6'h2d];
  assign T14162 = $signed(T14163) / $signed(22'h100000);
  assign T14163 = $signed(31'h457d965e) * $signed(16'h0);
  assign twiddle4_2_445_imag = T14168 + T14164;
  assign T14164 = {T14167, T14165};
  assign T14165 = $signed(T14166) / $signed(22'h100000);
  assign T14166 = $signed(30'h19937161) * $signed(16'hffff);
  assign T14167 = T14165[6'h2d:6'h2d];
  assign T14168 = $signed(T14169) / $signed(22'h100000);
  assign T14169 = $signed(31'h4555215b) * $signed(16'h0);
  assign T14170 = T10817[1'h0:1'h0];
  assign T14171 = T14184 ? twiddle4_2_447_imag : twiddle4_2_446_imag;
  assign twiddle4_2_446_imag = T14176 + T14172;
  assign T14172 = {T14175, T14173};
  assign T14173 = $signed(T14174) / $signed(22'h100000);
  assign T14174 = $signed(30'h19372a63) * $signed(16'hffff);
  assign T14175 = T14173[6'h2d:6'h2d];
  assign T14176 = $signed(T14177) / $signed(22'h100000);
  assign T14177 = $signed(31'h452d3d19) * $signed(16'h0);
  assign twiddle4_2_447_imag = T14182 + T14178;
  assign T14178 = {T14181, T14179};
  assign T14179 = $signed(T14180) / $signed(22'h100000);
  assign T14180 = $signed(30'h18daa52e) * $signed(16'hffff);
  assign T14181 = T14179[6'h2d:6'h2d];
  assign T14182 = $signed(T14183) / $signed(22'h100000);
  assign T14183 = $signed(31'h4505e9fb) * $signed(16'h0);
  assign T14184 = T10817[1'h0:1'h0];
  assign T14185 = T10817[1'h1:1'h1];
  assign T14186 = T10817[2'h2:2'h2];
  assign T14187 = T10817[2'h3:2'h3];
  assign T14188 = T10817[3'h4:3'h4];
  assign T14189 = T10817[3'h5:3'h5];
  assign T14190 = T14740 ? T14454 : T14191;
  assign T14191 = T14453 ? T14318 : T14192;
  assign T14192 = T14317 ? T14255 : T14193;
  assign T14193 = T14254 ? T14224 : T14194;
  assign T14194 = T14223 ? T14209 : T14195;
  assign T14195 = T14208 ? twiddle4_2_449_imag : twiddle4_2_448_imag;
  assign twiddle4_2_448_imag = T14200 + T14196;
  assign T14196 = {T14199, T14197};
  assign T14197 = $signed(T14198) / $signed(22'h100000);
  assign T14198 = $signed(30'h187de2a6) * $signed(16'hffff);
  assign T14199 = T14197[6'h2d:6'h2d];
  assign T14200 = $signed(T14201) / $signed(22'h100000);
  assign T14201 = $signed(31'h44df2862) * $signed(16'h0);
  assign twiddle4_2_449_imag = T14206 + T14202;
  assign T14202 = {T14205, T14203};
  assign T14203 = $signed(T14204) / $signed(22'h100000);
  assign T14204 = $signed(30'h1820e3b0) * $signed(16'hffff);
  assign T14205 = T14203[6'h2d:6'h2d];
  assign T14206 = $signed(T14207) / $signed(22'h100000);
  assign T14207 = $signed(31'h44b8f8ae) * $signed(16'h0);
  assign T14208 = T10817[1'h0:1'h0];
  assign T14209 = T14222 ? twiddle4_2_451_imag : twiddle4_2_450_imag;
  assign twiddle4_2_450_imag = T14214 + T14210;
  assign T14210 = {T14213, T14211};
  assign T14211 = $signed(T14212) / $signed(22'h100000);
  assign T14212 = $signed(30'h17c3a931) * $signed(16'hffff);
  assign T14213 = T14211[6'h2d:6'h2d];
  assign T14214 = $signed(T14215) / $signed(22'h100000);
  assign T14215 = $signed(31'h44935b3c) * $signed(16'h0);
  assign twiddle4_2_451_imag = T14220 + T14216;
  assign T14216 = {T14219, T14217};
  assign T14217 = $signed(T14218) / $signed(22'h100000);
  assign T14218 = $signed(30'h1766340f) * $signed(16'hffff);
  assign T14219 = T14217[6'h2d:6'h2d];
  assign T14220 = $signed(T14221) / $signed(22'h100000);
  assign T14221 = $signed(31'h446e506a) * $signed(16'h0);
  assign T14222 = T10817[1'h0:1'h0];
  assign T14223 = T10817[1'h1:1'h1];
  assign T14224 = T14253 ? T14239 : T14225;
  assign T14225 = T14238 ? twiddle4_2_453_imag : twiddle4_2_452_imag;
  assign twiddle4_2_452_imag = T14230 + T14226;
  assign T14226 = {T14229, T14227};
  assign T14227 = $signed(T14228) / $signed(22'h100000);
  assign T14228 = $signed(30'h17088530) * $signed(16'hffff);
  assign T14229 = T14227[6'h2d:6'h2d];
  assign T14230 = $signed(T14231) / $signed(22'h100000);
  assign T14231 = $signed(31'h4449d893) * $signed(16'h0);
  assign twiddle4_2_453_imag = T14236 + T14232;
  assign T14232 = {T14235, T14233};
  assign T14233 = $signed(T14234) / $signed(22'h100000);
  assign T14234 = $signed(30'h16aa9d7d) * $signed(16'hffff);
  assign T14235 = T14233[6'h2d:6'h2d];
  assign T14236 = $signed(T14237) / $signed(22'h100000);
  assign T14237 = $signed(31'h4425f411) * $signed(16'h0);
  assign T14238 = T10817[1'h0:1'h0];
  assign T14239 = T14252 ? twiddle4_2_455_imag : twiddle4_2_454_imag;
  assign twiddle4_2_454_imag = T14244 + T14240;
  assign T14240 = {T14243, T14241};
  assign T14241 = $signed(T14242) / $signed(22'h100000);
  assign T14242 = $signed(30'h164c7ddd) * $signed(16'hffff);
  assign T14243 = T14241[6'h2d:6'h2d];
  assign T14244 = $signed(T14245) / $signed(22'h100000);
  assign T14245 = $signed(31'h4402a33c) * $signed(16'h0);
  assign twiddle4_2_455_imag = T14250 + T14246;
  assign T14246 = {T14249, T14247};
  assign T14247 = $signed(T14248) / $signed(22'h100000);
  assign T14248 = $signed(30'h15ee2737) * $signed(16'hffff);
  assign T14249 = T14247[6'h2d:6'h2d];
  assign T14250 = $signed(T14251) / $signed(22'h100000);
  assign T14251 = $signed(31'h43dfe66c) * $signed(16'h0);
  assign T14252 = T10817[1'h0:1'h0];
  assign T14253 = T10817[1'h1:1'h1];
  assign T14254 = T10817[2'h2:2'h2];
  assign T14255 = T14316 ? T14286 : T14256;
  assign T14256 = T14285 ? T14271 : T14257;
  assign T14257 = T14270 ? twiddle4_2_457_imag : twiddle4_2_456_imag;
  assign twiddle4_2_456_imag = T14262 + T14258;
  assign T14258 = {T14261, T14259};
  assign T14259 = $signed(T14260) / $signed(22'h100000);
  assign T14260 = $signed(30'h158f9a75) * $signed(16'hffff);
  assign T14261 = T14259[6'h2d:6'h2d];
  assign T14262 = $signed(T14263) / $signed(22'h100000);
  assign T14263 = $signed(31'h43bdbdf7) * $signed(16'h0);
  assign twiddle4_2_457_imag = T14268 + T14264;
  assign T14264 = {T14267, T14265};
  assign T14265 = $signed(T14266) / $signed(22'h100000);
  assign T14266 = $signed(30'h1530d880) * $signed(16'hffff);
  assign T14267 = T14265[6'h2d:6'h2d];
  assign T14268 = $signed(T14269) / $signed(22'h100000);
  assign T14269 = $signed(31'h439c2a30) * $signed(16'h0);
  assign T14270 = T10817[1'h0:1'h0];
  assign T14271 = T14284 ? twiddle4_2_459_imag : twiddle4_2_458_imag;
  assign twiddle4_2_458_imag = T14276 + T14272;
  assign T14272 = {T14275, T14273};
  assign T14273 = $signed(T14274) / $signed(22'h100000);
  assign T14274 = $signed(30'h14d1e242) * $signed(16'hffff);
  assign T14275 = T14273[6'h2d:6'h2d];
  assign T14276 = $signed(T14277) / $signed(22'h100000);
  assign T14277 = $signed(31'h437b2b6a) * $signed(16'h0);
  assign twiddle4_2_459_imag = T14282 + T14278;
  assign T14278 = {T14281, T14279};
  assign T14279 = $signed(T14280) / $signed(22'h100000);
  assign T14280 = $signed(30'h1472b8a5) * $signed(16'hffff);
  assign T14281 = T14279[6'h2d:6'h2d];
  assign T14282 = $signed(T14283) / $signed(22'h100000);
  assign T14283 = $signed(31'h435ac1f8) * $signed(16'h0);
  assign T14284 = T10817[1'h0:1'h0];
  assign T14285 = T10817[1'h1:1'h1];
  assign T14286 = T14315 ? T14301 : T14287;
  assign T14287 = T14300 ? twiddle4_2_461_imag : twiddle4_2_460_imag;
  assign twiddle4_2_460_imag = T14292 + T14288;
  assign T14288 = {T14291, T14289};
  assign T14289 = $signed(T14290) / $signed(22'h100000);
  assign T14290 = $signed(30'h14135c94) * $signed(16'hffff);
  assign T14291 = T14289[6'h2d:6'h2d];
  assign T14292 = $signed(T14293) / $signed(22'h100000);
  assign T14293 = $signed(31'h433aee28) * $signed(16'h0);
  assign twiddle4_2_461_imag = T14298 + T14294;
  assign T14294 = {T14297, T14295};
  assign T14295 = $signed(T14296) / $signed(22'h100000);
  assign T14296 = $signed(30'h13b3cefa) * $signed(16'hffff);
  assign T14297 = T14295[6'h2d:6'h2d];
  assign T14298 = $signed(T14299) / $signed(22'h100000);
  assign T14299 = $signed(31'h431bb04a) * $signed(16'h0);
  assign T14300 = T10817[1'h0:1'h0];
  assign T14301 = T14314 ? twiddle4_2_463_imag : twiddle4_2_462_imag;
  assign twiddle4_2_462_imag = T14306 + T14302;
  assign T14302 = {T14305, T14303};
  assign T14303 = $signed(T14304) / $signed(22'h100000);
  assign T14304 = $signed(30'h135410c2) * $signed(16'hffff);
  assign T14305 = T14303[6'h2d:6'h2d];
  assign T14306 = $signed(T14307) / $signed(22'h100000);
  assign T14307 = $signed(31'h42fd08aa) * $signed(16'h0);
  assign twiddle4_2_463_imag = T14312 + T14308;
  assign T14308 = {T14311, T14309};
  assign T14309 = $signed(T14310) / $signed(22'h100000);
  assign T14310 = $signed(30'h12f422da) * $signed(16'hffff);
  assign T14311 = T14309[6'h2d:6'h2d];
  assign T14312 = $signed(T14313) / $signed(22'h100000);
  assign T14313 = $signed(31'h42def794) * $signed(16'h0);
  assign T14314 = T10817[1'h0:1'h0];
  assign T14315 = T10817[1'h1:1'h1];
  assign T14316 = T10817[2'h2:2'h2];
  assign T14317 = T10817[2'h3:2'h3];
  assign T14318 = T14452 ? T14382 : T14319;
  assign T14319 = T14381 ? T14350 : T14320;
  assign T14320 = T14349 ? T14335 : T14321;
  assign T14321 = T14334 ? twiddle4_2_465_imag : twiddle4_2_464_imag;
  assign twiddle4_2_464_imag = T14326 + T14322;
  assign T14322 = {T14325, T14323};
  assign T14323 = $signed(T14324) / $signed(22'h100000);
  assign T14324 = $signed(30'h1294062e) * $signed(16'hffff);
  assign T14325 = T14323[6'h2d:6'h2d];
  assign T14326 = $signed(T14327) / $signed(22'h100000);
  assign T14327 = $signed(31'h42c17d53) * $signed(16'h0);
  assign twiddle4_2_465_imag = T14332 + T14328;
  assign T14328 = {T14331, T14329};
  assign T14329 = $signed(T14330) / $signed(22'h100000);
  assign T14330 = $signed(30'h1233bbab) * $signed(16'hffff);
  assign T14331 = T14329[6'h2d:6'h2d];
  assign T14332 = $signed(T14333) / $signed(22'h100000);
  assign T14333 = $signed(31'h42a49a2f) * $signed(16'h0);
  assign T14334 = T10817[1'h0:1'h0];
  assign T14335 = T14348 ? twiddle4_2_467_imag : twiddle4_2_466_imag;
  assign twiddle4_2_466_imag = T14340 + T14336;
  assign T14336 = {T14339, T14337};
  assign T14337 = $signed(T14338) / $signed(22'h100000);
  assign T14338 = $signed(30'h11d3443f) * $signed(16'hffff);
  assign T14339 = T14337[6'h2d:6'h2d];
  assign T14340 = $signed(T14341) / $signed(22'h100000);
  assign T14341 = $signed(31'h42884e6f) * $signed(16'h0);
  assign twiddle4_2_467_imag = T14346 + T14342;
  assign T14342 = {T14345, T14343};
  assign T14343 = $signed(T14344) / $signed(22'h100000);
  assign T14344 = $signed(30'h1172a0d7) * $signed(16'hffff);
  assign T14345 = T14343[6'h2d:6'h2d];
  assign T14346 = $signed(T14347) / $signed(22'h100000);
  assign T14347 = $signed(31'h426c9a59) * $signed(16'h0);
  assign T14348 = T10817[1'h0:1'h0];
  assign T14349 = T10817[1'h1:1'h1];
  assign T14350 = T14380 ? T14365 : T14351;
  assign T14351 = T14364 ? twiddle4_2_469_imag : twiddle4_2_468_imag;
  assign twiddle4_2_468_imag = T14356 + T14352;
  assign T14352 = {T14355, T14353};
  assign T14353 = $signed(T14354) / $signed(22'h100000);
  assign T14354 = $signed(30'h1111d262) * $signed(16'hffff);
  assign T14355 = T14353[6'h2d:6'h2d];
  assign T14356 = $signed(T14357) / $signed(22'h100000);
  assign T14357 = $signed(31'h42517e32) * $signed(16'h0);
  assign twiddle4_2_469_imag = T14362 + T14358;
  assign T14358 = {T14361, T14359};
  assign T14359 = $signed(T14360) / $signed(22'h100000);
  assign T14360 = $signed(30'h10b0d9cf) * $signed(16'hffff);
  assign T14361 = T14359[6'h2d:6'h2d];
  assign T14362 = $signed(T14363) / $signed(22'h100000);
  assign T14363 = $signed(31'h4236fa3c) * $signed(16'h0);
  assign T14364 = T10817[1'h0:1'h0];
  assign T14365 = T14379 ? twiddle4_2_471_imag : twiddle4_2_470_imag;
  assign twiddle4_2_470_imag = T14370 + T14366;
  assign T14366 = {T14369, T14367};
  assign T14367 = $signed(T14368) / $signed(22'h100000);
  assign T14368 = $signed(30'h104fb80e) * $signed(16'hffff);
  assign T14369 = T14367[6'h2d:6'h2d];
  assign T14370 = $signed(T14371) / $signed(22'h100000);
  assign T14371 = $signed(31'h421d0eb9) * $signed(16'h0);
  assign twiddle4_2_471_imag = T14377 + T14372;
  assign T14372 = {T14375, T14373};
  assign T14373 = $signed(T14374) / $signed(22'h100000);
  assign T14374 = $signed(29'hfee6e0d) * $signed(16'hffff);
  assign T14375 = T14376 ? 2'h3 : 2'h0;
  assign T14376 = T14373[6'h2c:6'h2c];
  assign T14377 = $signed(T14378) / $signed(22'h100000);
  assign T14378 = $signed(31'h4203bbe8) * $signed(16'h0);
  assign T14379 = T10817[1'h0:1'h0];
  assign T14380 = T10817[1'h1:1'h1];
  assign T14381 = T10817[2'h2:2'h2];
  assign T14382 = T14451 ? T14417 : T14383;
  assign T14383 = T14416 ? T14400 : T14384;
  assign T14384 = T14399 ? twiddle4_2_473_imag : twiddle4_2_472_imag;
  assign twiddle4_2_472_imag = T14390 + T14385;
  assign T14385 = {T14388, T14386};
  assign T14386 = $signed(T14387) / $signed(22'h100000);
  assign T14387 = $signed(29'hf8cfcbd) * $signed(16'hffff);
  assign T14388 = T14389 ? 2'h3 : 2'h0;
  assign T14389 = T14386[6'h2c:6'h2c];
  assign T14390 = $signed(T14391) / $signed(22'h100000);
  assign T14391 = $signed(31'h41eb0209) * $signed(16'h0);
  assign twiddle4_2_473_imag = T14397 + T14392;
  assign T14392 = {T14395, T14393};
  assign T14393 = $signed(T14394) / $signed(22'h100000);
  assign T14394 = $signed(29'hf2b650f) * $signed(16'hffff);
  assign T14395 = T14396 ? 2'h3 : 2'h0;
  assign T14396 = T14393[6'h2c:6'h2c];
  assign T14397 = $signed(T14398) / $signed(22'h100000);
  assign T14398 = $signed(31'h41d2e159) * $signed(16'h0);
  assign T14399 = T10817[1'h0:1'h0];
  assign T14400 = T14415 ? twiddle4_2_475_imag : twiddle4_2_474_imag;
  assign twiddle4_2_474_imag = T14406 + T14401;
  assign T14401 = {T14404, T14402};
  assign T14402 = $signed(T14403) / $signed(22'h100000);
  assign T14403 = $signed(29'hec9a7f2) * $signed(16'hffff);
  assign T14404 = T14405 ? 2'h3 : 2'h0;
  assign T14405 = T14402[6'h2c:6'h2c];
  assign T14406 = $signed(T14407) / $signed(22'h100000);
  assign T14407 = $signed(31'h41bb5a12) * $signed(16'h0);
  assign twiddle4_2_475_imag = T14413 + T14408;
  assign T14408 = {T14411, T14409};
  assign T14409 = $signed(T14410) / $signed(22'h100000);
  assign T14410 = $signed(29'he67c659) * $signed(16'hffff);
  assign T14411 = T14412 ? 2'h3 : 2'h0;
  assign T14412 = T14409[6'h2c:6'h2c];
  assign T14413 = $signed(T14414) / $signed(22'h100000);
  assign T14414 = $signed(31'h41a46c6e) * $signed(16'h0);
  assign T14415 = T10817[1'h0:1'h0];
  assign T14416 = T10817[1'h1:1'h1];
  assign T14417 = T14450 ? T14434 : T14418;
  assign T14418 = T14433 ? twiddle4_2_477_imag : twiddle4_2_476_imag;
  assign twiddle4_2_476_imag = T14424 + T14419;
  assign T14419 = {T14422, T14420};
  assign T14420 = $signed(T14421) / $signed(22'h100000);
  assign T14421 = $signed(29'he05c135) * $signed(16'hffff);
  assign T14422 = T14423 ? 2'h3 : 2'h0;
  assign T14423 = T14420[6'h2c:6'h2c];
  assign T14424 = $signed(T14425) / $signed(22'h100000);
  assign T14425 = $signed(31'h418e18a8) * $signed(16'h0);
  assign twiddle4_2_477_imag = T14431 + T14426;
  assign T14426 = {T14429, T14427};
  assign T14427 = $signed(T14428) / $signed(22'h100000);
  assign T14428 = $signed(29'hda39977) * $signed(16'hffff);
  assign T14429 = T14430 ? 2'h3 : 2'h0;
  assign T14430 = T14427[6'h2c:6'h2c];
  assign T14431 = $signed(T14432) / $signed(22'h100000);
  assign T14432 = $signed(31'h41785ef5) * $signed(16'h0);
  assign T14433 = T10817[1'h0:1'h0];
  assign T14434 = T14449 ? twiddle4_2_479_imag : twiddle4_2_478_imag;
  assign twiddle4_2_478_imag = T14440 + T14435;
  assign T14435 = {T14438, T14436};
  assign T14436 = $signed(T14437) / $signed(22'h100000);
  assign T14437 = $signed(29'hd415012) * $signed(16'hffff);
  assign T14438 = T14439 ? 2'h3 : 2'h0;
  assign T14439 = T14436[6'h2c:6'h2c];
  assign T14440 = $signed(T14441) / $signed(22'h100000);
  assign T14441 = $signed(31'h41633f8a) * $signed(16'h0);
  assign twiddle4_2_479_imag = T14447 + T14442;
  assign T14442 = {T14445, T14443};
  assign T14443 = $signed(T14444) / $signed(22'h100000);
  assign T14444 = $signed(29'hcdee5f9) * $signed(16'hffff);
  assign T14445 = T14446 ? 2'h3 : 2'h0;
  assign T14446 = T14443[6'h2c:6'h2c];
  assign T14447 = $signed(T14448) / $signed(22'h100000);
  assign T14448 = $signed(31'h414eba9e) * $signed(16'h0);
  assign T14449 = T10817[1'h0:1'h0];
  assign T14450 = T10817[1'h1:1'h1];
  assign T14451 = T10817[2'h2:2'h2];
  assign T14452 = T10817[2'h3:2'h3];
  assign T14453 = T10817[3'h4:3'h4];
  assign T14454 = T14739 ? T14597 : T14455;
  assign T14455 = T14596 ? T14526 : T14456;
  assign T14456 = T14525 ? T14491 : T14457;
  assign T14457 = T14490 ? T14474 : T14458;
  assign T14458 = T14473 ? twiddle4_2_481_imag : twiddle4_2_480_imag;
  assign twiddle4_2_480_imag = T14464 + T14459;
  assign T14459 = {T14462, T14460};
  assign T14460 = $signed(T14461) / $signed(22'h100000);
  assign T14461 = $signed(29'hc7c5c1e) * $signed(16'hffff);
  assign T14462 = T14463 ? 2'h3 : 2'h0;
  assign T14463 = T14460[6'h2c:6'h2c];
  assign T14464 = $signed(T14465) / $signed(22'h100000);
  assign T14465 = $signed(31'h413ad061) * $signed(16'h0);
  assign twiddle4_2_481_imag = T14471 + T14466;
  assign T14466 = {T14469, T14467};
  assign T14467 = $signed(T14468) / $signed(22'h100000);
  assign T14468 = $signed(29'hc19b374) * $signed(16'hffff);
  assign T14469 = T14470 ? 2'h3 : 2'h0;
  assign T14470 = T14467[6'h2c:6'h2c];
  assign T14471 = $signed(T14472) / $signed(22'h100000);
  assign T14472 = $signed(31'h41278105) * $signed(16'h0);
  assign T14473 = T10817[1'h0:1'h0];
  assign T14474 = T14489 ? twiddle4_2_483_imag : twiddle4_2_482_imag;
  assign twiddle4_2_482_imag = T14480 + T14475;
  assign T14475 = {T14478, T14476};
  assign T14476 = $signed(T14477) / $signed(22'h100000);
  assign T14477 = $signed(29'hbb6ecef) * $signed(16'hffff);
  assign T14478 = T14479 ? 2'h3 : 2'h0;
  assign T14479 = T14476[6'h2c:6'h2c];
  assign T14480 = $signed(T14481) / $signed(22'h100000);
  assign T14481 = $signed(31'h4114ccb9) * $signed(16'h0);
  assign twiddle4_2_483_imag = T14487 + T14482;
  assign T14482 = {T14485, T14483};
  assign T14483 = $signed(T14484) / $signed(22'h100000);
  assign T14484 = $signed(29'hb540982) * $signed(16'hffff);
  assign T14485 = T14486 ? 2'h3 : 2'h0;
  assign T14486 = T14483[6'h2c:6'h2c];
  assign T14487 = $signed(T14488) / $signed(22'h100000);
  assign T14488 = $signed(31'h4102b3ad) * $signed(16'h0);
  assign T14489 = T10817[1'h0:1'h0];
  assign T14490 = T10817[1'h1:1'h1];
  assign T14491 = T14524 ? T14508 : T14492;
  assign T14492 = T14507 ? twiddle4_2_485_imag : twiddle4_2_484_imag;
  assign twiddle4_2_484_imag = T14498 + T14493;
  assign T14493 = {T14496, T14494};
  assign T14494 = $signed(T14495) / $signed(22'h100000);
  assign T14495 = $signed(29'haf10a22) * $signed(16'hffff);
  assign T14496 = T14497 ? 2'h3 : 2'h0;
  assign T14497 = T14494[6'h2c:6'h2c];
  assign T14498 = $signed(T14499) / $signed(22'h100000);
  assign T14499 = $signed(31'h40f1360c) * $signed(16'h0);
  assign twiddle4_2_485_imag = T14505 + T14500;
  assign T14500 = {T14503, T14501};
  assign T14501 = $signed(T14502) / $signed(22'h100000);
  assign T14502 = $signed(29'ha8defc2) * $signed(16'hffff);
  assign T14503 = T14504 ? 2'h3 : 2'h0;
  assign T14504 = T14501[6'h2c:6'h2c];
  assign T14505 = $signed(T14506) / $signed(22'h100000);
  assign T14506 = $signed(31'h40e05401) * $signed(16'h0);
  assign T14507 = T10817[1'h0:1'h0];
  assign T14508 = T14523 ? twiddle4_2_487_imag : twiddle4_2_486_imag;
  assign twiddle4_2_486_imag = T14514 + T14509;
  assign T14509 = {T14512, T14510};
  assign T14510 = $signed(T14511) / $signed(22'h100000);
  assign T14511 = $signed(29'ha2abb58) * $signed(16'hffff);
  assign T14512 = T14513 ? 2'h3 : 2'h0;
  assign T14513 = T14510[6'h2c:6'h2c];
  assign T14514 = $signed(T14515) / $signed(22'h100000);
  assign T14515 = $signed(31'h40d00db7) * $signed(16'h0);
  assign twiddle4_2_487_imag = T14521 + T14516;
  assign T14516 = {T14519, T14517};
  assign T14517 = $signed(T14518) / $signed(22'h100000);
  assign T14518 = $signed(29'h9c76dd8) * $signed(16'hffff);
  assign T14519 = T14520 ? 2'h3 : 2'h0;
  assign T14520 = T14517[6'h2c:6'h2c];
  assign T14521 = $signed(T14522) / $signed(22'h100000);
  assign T14522 = $signed(31'h40c06355) * $signed(16'h0);
  assign T14523 = T10817[1'h0:1'h0];
  assign T14524 = T10817[1'h1:1'h1];
  assign T14525 = T10817[2'h2:2'h2];
  assign T14526 = T14595 ? T14561 : T14527;
  assign T14527 = T14560 ? T14544 : T14528;
  assign T14528 = T14543 ? twiddle4_2_489_imag : twiddle4_2_488_imag;
  assign twiddle4_2_488_imag = T14534 + T14529;
  assign T14529 = {T14532, T14530};
  assign T14530 = $signed(T14531) / $signed(22'h100000);
  assign T14531 = $signed(29'h9640837) * $signed(16'hffff);
  assign T14532 = T14533 ? 2'h3 : 2'h0;
  assign T14533 = T14530[6'h2c:6'h2c];
  assign T14534 = $signed(T14535) / $signed(22'h100000);
  assign T14535 = $signed(31'h40b15502) * $signed(16'h0);
  assign twiddle4_2_489_imag = T14541 + T14536;
  assign T14536 = {T14539, T14537};
  assign T14537 = $signed(T14538) / $signed(22'h100000);
  assign T14538 = $signed(29'h9008b6a) * $signed(16'hffff);
  assign T14539 = T14540 ? 2'h3 : 2'h0;
  assign T14540 = T14537[6'h2c:6'h2c];
  assign T14541 = $signed(T14542) / $signed(22'h100000);
  assign T14542 = $signed(31'h40a2e2e4) * $signed(16'h0);
  assign T14543 = T10817[1'h0:1'h0];
  assign T14544 = T14559 ? twiddle4_2_491_imag : twiddle4_2_490_imag;
  assign twiddle4_2_490_imag = T14550 + T14545;
  assign T14545 = {T14548, T14546};
  assign T14546 = $signed(T14547) / $signed(22'h100000);
  assign T14547 = $signed(29'h89cf867) * $signed(16'hffff);
  assign T14548 = T14549 ? 2'h3 : 2'h0;
  assign T14549 = T14546[6'h2c:6'h2c];
  assign T14550 = $signed(T14551) / $signed(22'h100000);
  assign T14551 = $signed(31'h40950d1d) * $signed(16'h0);
  assign twiddle4_2_491_imag = T14557 + T14552;
  assign T14552 = {T14555, T14553};
  assign T14553 = $signed(T14554) / $signed(22'h100000);
  assign T14554 = $signed(29'h8395023) * $signed(16'hffff);
  assign T14555 = T14556 ? 2'h3 : 2'h0;
  assign T14556 = T14553[6'h2c:6'h2c];
  assign T14557 = $signed(T14558) / $signed(22'h100000);
  assign T14558 = $signed(31'h4087d3d1) * $signed(16'h0);
  assign T14559 = T10817[1'h0:1'h0];
  assign T14560 = T10817[1'h1:1'h1];
  assign T14561 = T14594 ? T14578 : T14562;
  assign T14562 = T14577 ? twiddle4_2_493_imag : twiddle4_2_492_imag;
  assign twiddle4_2_492_imag = T14568 + T14563;
  assign T14563 = {T14566, T14564};
  assign T14564 = $signed(T14565) / $signed(22'h100000);
  assign T14565 = $signed(28'h7d59395) * $signed(16'hffff);
  assign T14566 = T14567 ? 3'h7 : 3'h0;
  assign T14567 = T14564[6'h2b:6'h2b];
  assign T14568 = $signed(T14569) / $signed(22'h100000);
  assign T14569 = $signed(31'h407b371f) * $signed(16'h0);
  assign twiddle4_2_493_imag = T14575 + T14570;
  assign T14570 = {T14573, T14571};
  assign T14571 = $signed(T14572) / $signed(22'h100000);
  assign T14572 = $signed(28'h771c3b2) * $signed(16'hffff);
  assign T14573 = T14574 ? 3'h7 : 3'h0;
  assign T14574 = T14571[6'h2b:6'h2b];
  assign T14575 = $signed(T14576) / $signed(22'h100000);
  assign T14576 = $signed(31'h406f3727) * $signed(16'h0);
  assign T14577 = T10817[1'h0:1'h0];
  assign T14578 = T14593 ? twiddle4_2_495_imag : twiddle4_2_494_imag;
  assign twiddle4_2_494_imag = T14584 + T14579;
  assign T14579 = {T14582, T14580};
  assign T14580 = $signed(T14581) / $signed(22'h100000);
  assign T14581 = $signed(28'h70de171) * $signed(16'hffff);
  assign T14582 = T14583 ? 3'h7 : 3'h0;
  assign T14583 = T14580[6'h2b:6'h2b];
  assign T14584 = $signed(T14585) / $signed(22'h100000);
  assign T14585 = $signed(31'h4063d406) * $signed(16'h0);
  assign twiddle4_2_495_imag = T14591 + T14586;
  assign T14586 = {T14589, T14587};
  assign T14587 = $signed(T14588) / $signed(22'h100000);
  assign T14588 = $signed(28'h6a9edc9) * $signed(16'hffff);
  assign T14589 = T14590 ? 3'h7 : 3'h0;
  assign T14590 = T14587[6'h2b:6'h2b];
  assign T14591 = $signed(T14592) / $signed(22'h100000);
  assign T14592 = $signed(31'h40590dd8) * $signed(16'h0);
  assign T14593 = T10817[1'h0:1'h0];
  assign T14594 = T10817[1'h1:1'h1];
  assign T14595 = T10817[2'h2:2'h2];
  assign T14596 = T10817[2'h3:2'h3];
  assign T14597 = T14738 ? T14668 : T14598;
  assign T14598 = T14667 ? T14633 : T14599;
  assign T14599 = T14632 ? T14616 : T14600;
  assign T14600 = T14615 ? twiddle4_2_497_imag : twiddle4_2_496_imag;
  assign twiddle4_2_496_imag = T14606 + T14601;
  assign T14601 = {T14604, T14602};
  assign T14602 = $signed(T14603) / $signed(22'h100000);
  assign T14603 = $signed(28'h645e9af) * $signed(16'hffff);
  assign T14604 = T14605 ? 3'h7 : 3'h0;
  assign T14605 = T14602[6'h2b:6'h2b];
  assign T14606 = $signed(T14607) / $signed(22'h100000);
  assign T14607 = $signed(31'h404ee4b9) * $signed(16'h0);
  assign twiddle4_2_497_imag = T14613 + T14608;
  assign T14608 = {T14611, T14609};
  assign T14609 = $signed(T14610) / $signed(22'h100000);
  assign T14610 = $signed(28'h5e1d61a) * $signed(16'hffff);
  assign T14611 = T14612 ? 3'h7 : 3'h0;
  assign T14612 = T14609[6'h2b:6'h2b];
  assign T14613 = $signed(T14614) / $signed(22'h100000);
  assign T14614 = $signed(31'h404558c1) * $signed(16'h0);
  assign T14615 = T10817[1'h0:1'h0];
  assign T14616 = T14631 ? twiddle4_2_499_imag : twiddle4_2_498_imag;
  assign twiddle4_2_498_imag = T14622 + T14617;
  assign T14617 = {T14620, T14618};
  assign T14618 = $signed(T14619) / $signed(22'h100000);
  assign T14619 = $signed(28'h57db402) * $signed(16'hffff);
  assign T14620 = T14621 ? 3'h7 : 3'h0;
  assign T14621 = T14618[6'h2b:6'h2b];
  assign T14622 = $signed(T14623) / $signed(22'h100000);
  assign T14623 = $signed(31'h403c6a07) * $signed(16'h0);
  assign twiddle4_2_499_imag = T14629 + T14624;
  assign T14624 = {T14627, T14625};
  assign T14625 = $signed(T14626) / $signed(22'h100000);
  assign T14626 = $signed(28'h519845e) * $signed(16'hffff);
  assign T14627 = T14628 ? 3'h7 : 3'h0;
  assign T14628 = T14625[6'h2b:6'h2b];
  assign T14629 = $signed(T14630) / $signed(22'h100000);
  assign T14630 = $signed(31'h403418a2) * $signed(16'h0);
  assign T14631 = T10817[1'h0:1'h0];
  assign T14632 = T10817[1'h1:1'h1];
  assign T14633 = T14666 ? T14650 : T14634;
  assign T14634 = T14649 ? twiddle4_2_501_imag : twiddle4_2_500_imag;
  assign twiddle4_2_500_imag = T14640 + T14635;
  assign T14635 = {T14638, T14636};
  assign T14636 = $signed(T14637) / $signed(22'h100000);
  assign T14637 = $signed(28'h4b54824) * $signed(16'hffff);
  assign T14638 = T14639 ? 3'h7 : 3'h0;
  assign T14639 = T14636[6'h2b:6'h2b];
  assign T14640 = $signed(T14641) / $signed(22'h100000);
  assign T14641 = $signed(31'h402c64a6) * $signed(16'h0);
  assign twiddle4_2_501_imag = T14647 + T14642;
  assign T14642 = {T14645, T14643};
  assign T14643 = $signed(T14644) / $signed(22'h100000);
  assign T14644 = $signed(28'h451004d) * $signed(16'hffff);
  assign T14645 = T14646 ? 3'h7 : 3'h0;
  assign T14646 = T14643[6'h2b:6'h2b];
  assign T14647 = $signed(T14648) / $signed(22'h100000);
  assign T14648 = $signed(31'h40254e27) * $signed(16'h0);
  assign T14649 = T10817[1'h0:1'h0];
  assign T14650 = T14665 ? twiddle4_2_503_imag : twiddle4_2_502_imag;
  assign twiddle4_2_502_imag = T14656 + T14651;
  assign T14651 = {T14654, T14652};
  assign T14652 = $signed(T14653) / $signed(22'h100000);
  assign T14653 = $signed(27'h3ecadcf) * $signed(16'hffff);
  assign T14654 = T14655 ? 4'hf : 4'h0;
  assign T14655 = T14652[6'h2a:6'h2a];
  assign T14656 = $signed(T14657) / $signed(22'h100000);
  assign T14657 = $signed(31'h401ed535) * $signed(16'h0);
  assign twiddle4_2_503_imag = T14663 + T14658;
  assign T14658 = {T14661, T14659};
  assign T14659 = $signed(T14660) / $signed(22'h100000);
  assign T14660 = $signed(27'h38851a2) * $signed(16'hffff);
  assign T14661 = T14662 ? 4'hf : 4'h0;
  assign T14662 = T14659[6'h2a:6'h2a];
  assign T14663 = $signed(T14664) / $signed(22'h100000);
  assign T14664 = $signed(31'h4018f9e1) * $signed(16'h0);
  assign T14665 = T10817[1'h0:1'h0];
  assign T14666 = T10817[1'h1:1'h1];
  assign T14667 = T10817[2'h2:2'h2];
  assign T14668 = T14737 ? T14703 : T14669;
  assign T14669 = T14702 ? T14686 : T14670;
  assign T14670 = T14685 ? twiddle4_2_505_imag : twiddle4_2_504_imag;
  assign twiddle4_2_504_imag = T14676 + T14671;
  assign T14671 = {T14674, T14672};
  assign T14672 = $signed(T14673) / $signed(22'h100000);
  assign T14673 = $signed(27'h323ecbe) * $signed(16'hffff);
  assign T14674 = T14675 ? 4'hf : 4'h0;
  assign T14675 = T14672[6'h2a:6'h2a];
  assign T14676 = $signed(T14677) / $signed(22'h100000);
  assign T14677 = $signed(31'h4013bc3a) * $signed(16'h0);
  assign twiddle4_2_505_imag = T14683 + T14678;
  assign T14678 = {T14681, T14679};
  assign T14679 = $signed(T14680) / $signed(22'h100000);
  assign T14680 = $signed(27'h2bf801a) * $signed(16'hffff);
  assign T14681 = T14682 ? 4'hf : 4'h0;
  assign T14682 = T14679[6'h2a:6'h2a];
  assign T14683 = $signed(T14684) / $signed(22'h100000);
  assign T14684 = $signed(31'h400f1c4b) * $signed(16'h0);
  assign T14685 = T10817[1'h0:1'h0];
  assign T14686 = T14701 ? twiddle4_2_507_imag : twiddle4_2_506_imag;
  assign twiddle4_2_506_imag = T14692 + T14687;
  assign T14687 = {T14690, T14688};
  assign T14688 = $signed(T14689) / $signed(22'h100000);
  assign T14689 = $signed(27'h25b0cae) * $signed(16'hffff);
  assign T14690 = T14691 ? 4'hf : 4'h0;
  assign T14691 = T14688[6'h2a:6'h2a];
  assign T14692 = $signed(T14693) / $signed(22'h100000);
  assign T14693 = $signed(31'h400b1a21) * $signed(16'h0);
  assign twiddle4_2_507_imag = T14699 + T14694;
  assign T14694 = {T14697, T14695};
  assign T14695 = $signed(T14696) / $signed(22'h100000);
  assign T14696 = $signed(26'h1f69373) * $signed(16'hffff);
  assign T14697 = T14698 ? 5'h1f : 5'h0;
  assign T14698 = T14695[6'h29:6'h29];
  assign T14699 = $signed(T14700) / $signed(22'h100000);
  assign T14700 = $signed(31'h4007b5c5) * $signed(16'h0);
  assign T14701 = T10817[1'h0:1'h0];
  assign T14702 = T10817[1'h1:1'h1];
  assign T14703 = T14736 ? T14720 : T14704;
  assign T14704 = T14719 ? twiddle4_2_509_imag : twiddle4_2_508_imag;
  assign twiddle4_2_508_imag = T14710 + T14705;
  assign T14705 = {T14708, T14706};
  assign T14706 = $signed(T14707) / $signed(22'h100000);
  assign T14707 = $signed(26'h192155f) * $signed(16'hffff);
  assign T14708 = T14709 ? 5'h1f : 5'h0;
  assign T14709 = T14706[6'h29:6'h29];
  assign T14710 = $signed(T14711) / $signed(22'h100000);
  assign T14711 = $signed(31'h4004ef3f) * $signed(16'h0);
  assign twiddle4_2_509_imag = T14717 + T14712;
  assign T14712 = {T14715, T14713};
  assign T14713 = $signed(T14714) / $signed(22'h100000);
  assign T14714 = $signed(26'h12d936b) * $signed(16'hffff);
  assign T14715 = T14716 ? 5'h1f : 5'h0;
  assign T14716 = T14713[6'h29:6'h29];
  assign T14717 = $signed(T14718) / $signed(22'h100000);
  assign T14718 = $signed(31'h4002c698) * $signed(16'h0);
  assign T14719 = T10817[1'h0:1'h0];
  assign T14720 = T14735 ? twiddle4_2_511_imag : twiddle4_2_510_imag;
  assign twiddle4_2_510_imag = T14726 + T14721;
  assign T14721 = {T14724, T14722};
  assign T14722 = $signed(T14723) / $signed(22'h100000);
  assign T14723 = $signed(25'hc90e8f) * $signed(16'hffff);
  assign T14724 = T14725 ? 6'h3f : 6'h0;
  assign T14725 = T14722[6'h28:6'h28];
  assign T14726 = $signed(T14727) / $signed(22'h100000);
  assign T14727 = $signed(31'h40013bd3) * $signed(16'h0);
  assign twiddle4_2_511_imag = T14733 + T14728;
  assign T14728 = {T14731, T14729};
  assign T14729 = $signed(T14730) / $signed(22'h100000);
  assign T14730 = $signed(24'h6487c3) * $signed(16'hffff);
  assign T14731 = T14732 ? 7'h7f : 7'h0;
  assign T14732 = T14729[6'h27:6'h27];
  assign T14733 = $signed(T14734) / $signed(22'h100000);
  assign T14734 = $signed(31'h40004ef5) * $signed(16'h0);
  assign T14735 = T10817[1'h0:1'h0];
  assign T14736 = T10817[1'h1:1'h1];
  assign T14737 = T10817[2'h2:2'h2];
  assign T14738 = T10817[2'h3:2'h3];
  assign T14739 = T10817[3'h4:3'h4];
  assign T14740 = T10817[3'h5:3'h5];
  assign T14741 = T10817[3'h6:3'h6];
  assign T14742 = T13765[6'h2e:6'h2e];
  assign T14743 = T10817[3'h7:3'h7];
  assign T14744 = T10817[4'h8:4'h8];
  assign io_t4_2out_real = T14745;
  assign T14745 = T14746[4'hf:1'h0];
  assign T14746 = T18697 ? T16722 : T14747;
  assign T14747 = T16721 ? T15742 : T14748;
  assign T14748 = T15741 ? T15313 : T14749;
  assign T14749 = T15312 ? T15046 : T14750;
  assign T14750 = T15045 ? T14901 : T14751;
  assign T14751 = T14900 ? T14828 : T14752;
  assign T14752 = T14827 ? T14791 : T14753;
  assign T14753 = T14790 ? T14772 : T14754;
  assign T14754 = T14771 ? T14762 : twiddle4_2_0_real;
  assign twiddle4_2_0_real = T14760 + T14755;
  assign T14755 = {T14758, T14756};
  assign T14756 = $signed(T14757) / $signed(22'h100000);
  assign T14757 = $signed(1'h0) * $signed(16'h0);
  assign T14758 = T14759 ? 31'h7fffffff : 31'h0;
  assign T14759 = T14756[5'h10:5'h10];
  assign T14760 = $signed(T14761) / $signed(22'h100000);
  assign T14761 = $signed(32'h40000000) * $signed(16'h1);
  assign T14762 = {T14770, twiddle4_2_1_real};
  assign twiddle4_2_1_real = T14768 + T14763;
  assign T14763 = {T14766, T14764};
  assign T14764 = $signed(T14765) / $signed(22'h100000);
  assign T14765 = $signed(24'h6487c3) * $signed(16'h0);
  assign T14766 = T14767 ? 7'h7f : 7'h0;
  assign T14767 = T14764[6'h27:6'h27];
  assign T14768 = $signed(T14769) / $signed(22'h100000);
  assign T14769 = $signed(31'h3fffb10b) * $signed(16'h1);
  assign T14770 = twiddle4_2_1_real[6'h2e:6'h2e];
  assign T14771 = T10817[1'h0:1'h0];
  assign T14772 = {T14789, T14773};
  assign T14773 = T14788 ? twiddle4_2_3_real : twiddle4_2_2_real;
  assign twiddle4_2_2_real = T14779 + T14774;
  assign T14774 = {T14777, T14775};
  assign T14775 = $signed(T14776) / $signed(22'h100000);
  assign T14776 = $signed(25'hc90e8f) * $signed(16'h0);
  assign T14777 = T14778 ? 6'h3f : 6'h0;
  assign T14778 = T14775[6'h28:6'h28];
  assign T14779 = $signed(T14780) / $signed(22'h100000);
  assign T14780 = $signed(31'h3ffec42d) * $signed(16'h1);
  assign twiddle4_2_3_real = T14786 + T14781;
  assign T14781 = {T14784, T14782};
  assign T14782 = $signed(T14783) / $signed(22'h100000);
  assign T14783 = $signed(26'h12d936b) * $signed(16'h0);
  assign T14784 = T14785 ? 5'h1f : 5'h0;
  assign T14785 = T14782[6'h29:6'h29];
  assign T14786 = $signed(T14787) / $signed(22'h100000);
  assign T14787 = $signed(31'h3ffd3968) * $signed(16'h1);
  assign T14788 = T10817[1'h0:1'h0];
  assign T14789 = T14773[6'h2e:6'h2e];
  assign T14790 = T10817[1'h1:1'h1];
  assign T14791 = {T14826, T14792};
  assign T14792 = T14825 ? T14809 : T14793;
  assign T14793 = T14808 ? twiddle4_2_5_real : twiddle4_2_4_real;
  assign twiddle4_2_4_real = T14799 + T14794;
  assign T14794 = {T14797, T14795};
  assign T14795 = $signed(T14796) / $signed(22'h100000);
  assign T14796 = $signed(26'h192155f) * $signed(16'h0);
  assign T14797 = T14798 ? 5'h1f : 5'h0;
  assign T14798 = T14795[6'h29:6'h29];
  assign T14799 = $signed(T14800) / $signed(22'h100000);
  assign T14800 = $signed(31'h3ffb10c1) * $signed(16'h1);
  assign twiddle4_2_5_real = T14806 + T14801;
  assign T14801 = {T14804, T14802};
  assign T14802 = $signed(T14803) / $signed(22'h100000);
  assign T14803 = $signed(26'h1f69373) * $signed(16'h0);
  assign T14804 = T14805 ? 5'h1f : 5'h0;
  assign T14805 = T14802[6'h29:6'h29];
  assign T14806 = $signed(T14807) / $signed(22'h100000);
  assign T14807 = $signed(31'h3ff84a3b) * $signed(16'h1);
  assign T14808 = T10817[1'h0:1'h0];
  assign T14809 = T14824 ? twiddle4_2_7_real : twiddle4_2_6_real;
  assign twiddle4_2_6_real = T14815 + T14810;
  assign T14810 = {T14813, T14811};
  assign T14811 = $signed(T14812) / $signed(22'h100000);
  assign T14812 = $signed(27'h25b0cae) * $signed(16'h0);
  assign T14813 = T14814 ? 4'hf : 4'h0;
  assign T14814 = T14811[6'h2a:6'h2a];
  assign T14815 = $signed(T14816) / $signed(22'h100000);
  assign T14816 = $signed(31'h3ff4e5df) * $signed(16'h1);
  assign twiddle4_2_7_real = T14822 + T14817;
  assign T14817 = {T14820, T14818};
  assign T14818 = $signed(T14819) / $signed(22'h100000);
  assign T14819 = $signed(27'h2bf801a) * $signed(16'h0);
  assign T14820 = T14821 ? 4'hf : 4'h0;
  assign T14821 = T14818[6'h2a:6'h2a];
  assign T14822 = $signed(T14823) / $signed(22'h100000);
  assign T14823 = $signed(31'h3ff0e3b5) * $signed(16'h1);
  assign T14824 = T10817[1'h0:1'h0];
  assign T14825 = T10817[1'h1:1'h1];
  assign T14826 = T14792[6'h2e:6'h2e];
  assign T14827 = T10817[2'h2:2'h2];
  assign T14828 = {T14899, T14829};
  assign T14829 = T14898 ? T14864 : T14830;
  assign T14830 = T14863 ? T14847 : T14831;
  assign T14831 = T14846 ? twiddle4_2_9_real : twiddle4_2_8_real;
  assign twiddle4_2_8_real = T14837 + T14832;
  assign T14832 = {T14835, T14833};
  assign T14833 = $signed(T14834) / $signed(22'h100000);
  assign T14834 = $signed(27'h323ecbe) * $signed(16'h0);
  assign T14835 = T14836 ? 4'hf : 4'h0;
  assign T14836 = T14833[6'h2a:6'h2a];
  assign T14837 = $signed(T14838) / $signed(22'h100000);
  assign T14838 = $signed(31'h3fec43c6) * $signed(16'h1);
  assign twiddle4_2_9_real = T14844 + T14839;
  assign T14839 = {T14842, T14840};
  assign T14840 = $signed(T14841) / $signed(22'h100000);
  assign T14841 = $signed(27'h38851a2) * $signed(16'h0);
  assign T14842 = T14843 ? 4'hf : 4'h0;
  assign T14843 = T14840[6'h2a:6'h2a];
  assign T14844 = $signed(T14845) / $signed(22'h100000);
  assign T14845 = $signed(31'h3fe7061f) * $signed(16'h1);
  assign T14846 = T10817[1'h0:1'h0];
  assign T14847 = T14862 ? twiddle4_2_11_real : twiddle4_2_10_real;
  assign twiddle4_2_10_real = T14853 + T14848;
  assign T14848 = {T14851, T14849};
  assign T14849 = $signed(T14850) / $signed(22'h100000);
  assign T14850 = $signed(27'h3ecadcf) * $signed(16'h0);
  assign T14851 = T14852 ? 4'hf : 4'h0;
  assign T14852 = T14849[6'h2a:6'h2a];
  assign T14853 = $signed(T14854) / $signed(22'h100000);
  assign T14854 = $signed(31'h3fe12acb) * $signed(16'h1);
  assign twiddle4_2_11_real = T14860 + T14855;
  assign T14855 = {T14858, T14856};
  assign T14856 = $signed(T14857) / $signed(22'h100000);
  assign T14857 = $signed(28'h451004d) * $signed(16'h0);
  assign T14858 = T14859 ? 3'h7 : 3'h0;
  assign T14859 = T14856[6'h2b:6'h2b];
  assign T14860 = $signed(T14861) / $signed(22'h100000);
  assign T14861 = $signed(31'h3fdab1d9) * $signed(16'h1);
  assign T14862 = T10817[1'h0:1'h0];
  assign T14863 = T10817[1'h1:1'h1];
  assign T14864 = T14897 ? T14881 : T14865;
  assign T14865 = T14880 ? twiddle4_2_13_real : twiddle4_2_12_real;
  assign twiddle4_2_12_real = T14871 + T14866;
  assign T14866 = {T14869, T14867};
  assign T14867 = $signed(T14868) / $signed(22'h100000);
  assign T14868 = $signed(28'h4b54824) * $signed(16'h0);
  assign T14869 = T14870 ? 3'h7 : 3'h0;
  assign T14870 = T14867[6'h2b:6'h2b];
  assign T14871 = $signed(T14872) / $signed(22'h100000);
  assign T14872 = $signed(31'h3fd39b5a) * $signed(16'h1);
  assign twiddle4_2_13_real = T14878 + T14873;
  assign T14873 = {T14876, T14874};
  assign T14874 = $signed(T14875) / $signed(22'h100000);
  assign T14875 = $signed(28'h519845e) * $signed(16'h0);
  assign T14876 = T14877 ? 3'h7 : 3'h0;
  assign T14877 = T14874[6'h2b:6'h2b];
  assign T14878 = $signed(T14879) / $signed(22'h100000);
  assign T14879 = $signed(31'h3fcbe75e) * $signed(16'h1);
  assign T14880 = T10817[1'h0:1'h0];
  assign T14881 = T14896 ? twiddle4_2_15_real : twiddle4_2_14_real;
  assign twiddle4_2_14_real = T14887 + T14882;
  assign T14882 = {T14885, T14883};
  assign T14883 = $signed(T14884) / $signed(22'h100000);
  assign T14884 = $signed(28'h57db402) * $signed(16'h0);
  assign T14885 = T14886 ? 3'h7 : 3'h0;
  assign T14886 = T14883[6'h2b:6'h2b];
  assign T14887 = $signed(T14888) / $signed(22'h100000);
  assign T14888 = $signed(31'h3fc395f9) * $signed(16'h1);
  assign twiddle4_2_15_real = T14894 + T14889;
  assign T14889 = {T14892, T14890};
  assign T14890 = $signed(T14891) / $signed(22'h100000);
  assign T14891 = $signed(28'h5e1d61a) * $signed(16'h0);
  assign T14892 = T14893 ? 3'h7 : 3'h0;
  assign T14893 = T14890[6'h2b:6'h2b];
  assign T14894 = $signed(T14895) / $signed(22'h100000);
  assign T14895 = $signed(31'h3fbaa73f) * $signed(16'h1);
  assign T14896 = T10817[1'h0:1'h0];
  assign T14897 = T10817[1'h1:1'h1];
  assign T14898 = T10817[2'h2:2'h2];
  assign T14899 = T14829[6'h2e:6'h2e];
  assign T14900 = T10817[2'h3:2'h3];
  assign T14901 = {T15044, T14902};
  assign T14902 = T15043 ? T14973 : T14903;
  assign T14903 = T14972 ? T14938 : T14904;
  assign T14904 = T14937 ? T14921 : T14905;
  assign T14905 = T14920 ? twiddle4_2_17_real : twiddle4_2_16_real;
  assign twiddle4_2_16_real = T14911 + T14906;
  assign T14906 = {T14909, T14907};
  assign T14907 = $signed(T14908) / $signed(22'h100000);
  assign T14908 = $signed(28'h645e9af) * $signed(16'h0);
  assign T14909 = T14910 ? 3'h7 : 3'h0;
  assign T14910 = T14907[6'h2b:6'h2b];
  assign T14911 = $signed(T14912) / $signed(22'h100000);
  assign T14912 = $signed(31'h3fb11b47) * $signed(16'h1);
  assign twiddle4_2_17_real = T14918 + T14913;
  assign T14913 = {T14916, T14914};
  assign T14914 = $signed(T14915) / $signed(22'h100000);
  assign T14915 = $signed(28'h6a9edc9) * $signed(16'h0);
  assign T14916 = T14917 ? 3'h7 : 3'h0;
  assign T14917 = T14914[6'h2b:6'h2b];
  assign T14918 = $signed(T14919) / $signed(22'h100000);
  assign T14919 = $signed(31'h3fa6f228) * $signed(16'h1);
  assign T14920 = T10817[1'h0:1'h0];
  assign T14921 = T14936 ? twiddle4_2_19_real : twiddle4_2_18_real;
  assign twiddle4_2_18_real = T14927 + T14922;
  assign T14922 = {T14925, T14923};
  assign T14923 = $signed(T14924) / $signed(22'h100000);
  assign T14924 = $signed(28'h70de171) * $signed(16'h0);
  assign T14925 = T14926 ? 3'h7 : 3'h0;
  assign T14926 = T14923[6'h2b:6'h2b];
  assign T14927 = $signed(T14928) / $signed(22'h100000);
  assign T14928 = $signed(31'h3f9c2bfa) * $signed(16'h1);
  assign twiddle4_2_19_real = T14934 + T14929;
  assign T14929 = {T14932, T14930};
  assign T14930 = $signed(T14931) / $signed(22'h100000);
  assign T14931 = $signed(28'h771c3b2) * $signed(16'h0);
  assign T14932 = T14933 ? 3'h7 : 3'h0;
  assign T14933 = T14930[6'h2b:6'h2b];
  assign T14934 = $signed(T14935) / $signed(22'h100000);
  assign T14935 = $signed(31'h3f90c8d9) * $signed(16'h1);
  assign T14936 = T10817[1'h0:1'h0];
  assign T14937 = T10817[1'h1:1'h1];
  assign T14938 = T14971 ? T14955 : T14939;
  assign T14939 = T14954 ? twiddle4_2_21_real : twiddle4_2_20_real;
  assign twiddle4_2_20_real = T14945 + T14940;
  assign T14940 = {T14943, T14941};
  assign T14941 = $signed(T14942) / $signed(22'h100000);
  assign T14942 = $signed(28'h7d59395) * $signed(16'h0);
  assign T14943 = T14944 ? 3'h7 : 3'h0;
  assign T14944 = T14941[6'h2b:6'h2b];
  assign T14945 = $signed(T14946) / $signed(22'h100000);
  assign T14946 = $signed(31'h3f84c8e1) * $signed(16'h1);
  assign twiddle4_2_21_real = T14952 + T14947;
  assign T14947 = {T14950, T14948};
  assign T14948 = $signed(T14949) / $signed(22'h100000);
  assign T14949 = $signed(29'h8395023) * $signed(16'h0);
  assign T14950 = T14951 ? 2'h3 : 2'h0;
  assign T14951 = T14948[6'h2c:6'h2c];
  assign T14952 = $signed(T14953) / $signed(22'h100000);
  assign T14953 = $signed(31'h3f782c2f) * $signed(16'h1);
  assign T14954 = T10817[1'h0:1'h0];
  assign T14955 = T14970 ? twiddle4_2_23_real : twiddle4_2_22_real;
  assign twiddle4_2_22_real = T14961 + T14956;
  assign T14956 = {T14959, T14957};
  assign T14957 = $signed(T14958) / $signed(22'h100000);
  assign T14958 = $signed(29'h89cf867) * $signed(16'h0);
  assign T14959 = T14960 ? 2'h3 : 2'h0;
  assign T14960 = T14957[6'h2c:6'h2c];
  assign T14961 = $signed(T14962) / $signed(22'h100000);
  assign T14962 = $signed(31'h3f6af2e3) * $signed(16'h1);
  assign twiddle4_2_23_real = T14968 + T14963;
  assign T14963 = {T14966, T14964};
  assign T14964 = $signed(T14965) / $signed(22'h100000);
  assign T14965 = $signed(29'h9008b6a) * $signed(16'h0);
  assign T14966 = T14967 ? 2'h3 : 2'h0;
  assign T14967 = T14964[6'h2c:6'h2c];
  assign T14968 = $signed(T14969) / $signed(22'h100000);
  assign T14969 = $signed(31'h3f5d1d1c) * $signed(16'h1);
  assign T14970 = T10817[1'h0:1'h0];
  assign T14971 = T10817[1'h1:1'h1];
  assign T14972 = T10817[2'h2:2'h2];
  assign T14973 = T15042 ? T15008 : T14974;
  assign T14974 = T15007 ? T14991 : T14975;
  assign T14975 = T14990 ? twiddle4_2_25_real : twiddle4_2_24_real;
  assign twiddle4_2_24_real = T14981 + T14976;
  assign T14976 = {T14979, T14977};
  assign T14977 = $signed(T14978) / $signed(22'h100000);
  assign T14978 = $signed(29'h9640837) * $signed(16'h0);
  assign T14979 = T14980 ? 2'h3 : 2'h0;
  assign T14980 = T14977[6'h2c:6'h2c];
  assign T14981 = $signed(T14982) / $signed(22'h100000);
  assign T14982 = $signed(31'h3f4eaafe) * $signed(16'h1);
  assign twiddle4_2_25_real = T14988 + T14983;
  assign T14983 = {T14986, T14984};
  assign T14984 = $signed(T14985) / $signed(22'h100000);
  assign T14985 = $signed(29'h9c76dd8) * $signed(16'h0);
  assign T14986 = T14987 ? 2'h3 : 2'h0;
  assign T14987 = T14984[6'h2c:6'h2c];
  assign T14988 = $signed(T14989) / $signed(22'h100000);
  assign T14989 = $signed(31'h3f3f9cab) * $signed(16'h1);
  assign T14990 = T10817[1'h0:1'h0];
  assign T14991 = T15006 ? twiddle4_2_27_real : twiddle4_2_26_real;
  assign twiddle4_2_26_real = T14997 + T14992;
  assign T14992 = {T14995, T14993};
  assign T14993 = $signed(T14994) / $signed(22'h100000);
  assign T14994 = $signed(29'ha2abb58) * $signed(16'h0);
  assign T14995 = T14996 ? 2'h3 : 2'h0;
  assign T14996 = T14993[6'h2c:6'h2c];
  assign T14997 = $signed(T14998) / $signed(22'h100000);
  assign T14998 = $signed(31'h3f2ff249) * $signed(16'h1);
  assign twiddle4_2_27_real = T15004 + T14999;
  assign T14999 = {T15002, T15000};
  assign T15000 = $signed(T15001) / $signed(22'h100000);
  assign T15001 = $signed(29'ha8defc2) * $signed(16'h0);
  assign T15002 = T15003 ? 2'h3 : 2'h0;
  assign T15003 = T15000[6'h2c:6'h2c];
  assign T15004 = $signed(T15005) / $signed(22'h100000);
  assign T15005 = $signed(31'h3f1fabff) * $signed(16'h1);
  assign T15006 = T10817[1'h0:1'h0];
  assign T15007 = T10817[1'h1:1'h1];
  assign T15008 = T15041 ? T15025 : T15009;
  assign T15009 = T15024 ? twiddle4_2_29_real : twiddle4_2_28_real;
  assign twiddle4_2_28_real = T15015 + T15010;
  assign T15010 = {T15013, T15011};
  assign T15011 = $signed(T15012) / $signed(22'h100000);
  assign T15012 = $signed(29'haf10a22) * $signed(16'h0);
  assign T15013 = T15014 ? 2'h3 : 2'h0;
  assign T15014 = T15011[6'h2c:6'h2c];
  assign T15015 = $signed(T15016) / $signed(22'h100000);
  assign T15016 = $signed(31'h3f0ec9f4) * $signed(16'h1);
  assign twiddle4_2_29_real = T15022 + T15017;
  assign T15017 = {T15020, T15018};
  assign T15018 = $signed(T15019) / $signed(22'h100000);
  assign T15019 = $signed(29'hb540982) * $signed(16'h0);
  assign T15020 = T15021 ? 2'h3 : 2'h0;
  assign T15021 = T15018[6'h2c:6'h2c];
  assign T15022 = $signed(T15023) / $signed(22'h100000);
  assign T15023 = $signed(31'h3efd4c53) * $signed(16'h1);
  assign T15024 = T10817[1'h0:1'h0];
  assign T15025 = T15040 ? twiddle4_2_31_real : twiddle4_2_30_real;
  assign twiddle4_2_30_real = T15031 + T15026;
  assign T15026 = {T15029, T15027};
  assign T15027 = $signed(T15028) / $signed(22'h100000);
  assign T15028 = $signed(29'hbb6ecef) * $signed(16'h0);
  assign T15029 = T15030 ? 2'h3 : 2'h0;
  assign T15030 = T15027[6'h2c:6'h2c];
  assign T15031 = $signed(T15032) / $signed(22'h100000);
  assign T15032 = $signed(31'h3eeb3347) * $signed(16'h1);
  assign twiddle4_2_31_real = T15038 + T15033;
  assign T15033 = {T15036, T15034};
  assign T15034 = $signed(T15035) / $signed(22'h100000);
  assign T15035 = $signed(29'hc19b374) * $signed(16'h0);
  assign T15036 = T15037 ? 2'h3 : 2'h0;
  assign T15037 = T15034[6'h2c:6'h2c];
  assign T15038 = $signed(T15039) / $signed(22'h100000);
  assign T15039 = $signed(31'h3ed87efb) * $signed(16'h1);
  assign T15040 = T10817[1'h0:1'h0];
  assign T15041 = T10817[1'h1:1'h1];
  assign T15042 = T10817[2'h2:2'h2];
  assign T15043 = T10817[2'h3:2'h3];
  assign T15044 = T14902[6'h2e:6'h2e];
  assign T15045 = T10817[3'h4:3'h4];
  assign T15046 = {T15311, T15047};
  assign T15047 = T15310 ? T15184 : T15048;
  assign T15048 = T15183 ? T15119 : T15049;
  assign T15049 = T15118 ? T15084 : T15050;
  assign T15050 = T15083 ? T15067 : T15051;
  assign T15051 = T15066 ? twiddle4_2_33_real : twiddle4_2_32_real;
  assign twiddle4_2_32_real = T15057 + T15052;
  assign T15052 = {T15055, T15053};
  assign T15053 = $signed(T15054) / $signed(22'h100000);
  assign T15054 = $signed(29'hc7c5c1e) * $signed(16'h0);
  assign T15055 = T15056 ? 2'h3 : 2'h0;
  assign T15056 = T15053[6'h2c:6'h2c];
  assign T15057 = $signed(T15058) / $signed(22'h100000);
  assign T15058 = $signed(31'h3ec52f9f) * $signed(16'h1);
  assign twiddle4_2_33_real = T15064 + T15059;
  assign T15059 = {T15062, T15060};
  assign T15060 = $signed(T15061) / $signed(22'h100000);
  assign T15061 = $signed(29'hcdee5f9) * $signed(16'h0);
  assign T15062 = T15063 ? 2'h3 : 2'h0;
  assign T15063 = T15060[6'h2c:6'h2c];
  assign T15064 = $signed(T15065) / $signed(22'h100000);
  assign T15065 = $signed(31'h3eb14562) * $signed(16'h1);
  assign T15066 = T10817[1'h0:1'h0];
  assign T15067 = T15082 ? twiddle4_2_35_real : twiddle4_2_34_real;
  assign twiddle4_2_34_real = T15073 + T15068;
  assign T15068 = {T15071, T15069};
  assign T15069 = $signed(T15070) / $signed(22'h100000);
  assign T15070 = $signed(29'hd415012) * $signed(16'h0);
  assign T15071 = T15072 ? 2'h3 : 2'h0;
  assign T15072 = T15069[6'h2c:6'h2c];
  assign T15073 = $signed(T15074) / $signed(22'h100000);
  assign T15074 = $signed(31'h3e9cc076) * $signed(16'h1);
  assign twiddle4_2_35_real = T15080 + T15075;
  assign T15075 = {T15078, T15076};
  assign T15076 = $signed(T15077) / $signed(22'h100000);
  assign T15077 = $signed(29'hda39977) * $signed(16'h0);
  assign T15078 = T15079 ? 2'h3 : 2'h0;
  assign T15079 = T15076[6'h2c:6'h2c];
  assign T15080 = $signed(T15081) / $signed(22'h100000);
  assign T15081 = $signed(31'h3e87a10b) * $signed(16'h1);
  assign T15082 = T10817[1'h0:1'h0];
  assign T15083 = T10817[1'h1:1'h1];
  assign T15084 = T15117 ? T15101 : T15085;
  assign T15085 = T15100 ? twiddle4_2_37_real : twiddle4_2_36_real;
  assign twiddle4_2_36_real = T15091 + T15086;
  assign T15086 = {T15089, T15087};
  assign T15087 = $signed(T15088) / $signed(22'h100000);
  assign T15088 = $signed(29'he05c135) * $signed(16'h0);
  assign T15089 = T15090 ? 2'h3 : 2'h0;
  assign T15090 = T15087[6'h2c:6'h2c];
  assign T15091 = $signed(T15092) / $signed(22'h100000);
  assign T15092 = $signed(31'h3e71e758) * $signed(16'h1);
  assign twiddle4_2_37_real = T15098 + T15093;
  assign T15093 = {T15096, T15094};
  assign T15094 = $signed(T15095) / $signed(22'h100000);
  assign T15095 = $signed(29'he67c659) * $signed(16'h0);
  assign T15096 = T15097 ? 2'h3 : 2'h0;
  assign T15097 = T15094[6'h2c:6'h2c];
  assign T15098 = $signed(T15099) / $signed(22'h100000);
  assign T15099 = $signed(31'h3e5b9392) * $signed(16'h1);
  assign T15100 = T10817[1'h0:1'h0];
  assign T15101 = T15116 ? twiddle4_2_39_real : twiddle4_2_38_real;
  assign twiddle4_2_38_real = T15107 + T15102;
  assign T15102 = {T15105, T15103};
  assign T15103 = $signed(T15104) / $signed(22'h100000);
  assign T15104 = $signed(29'hec9a7f2) * $signed(16'h0);
  assign T15105 = T15106 ? 2'h3 : 2'h0;
  assign T15106 = T15103[6'h2c:6'h2c];
  assign T15107 = $signed(T15108) / $signed(22'h100000);
  assign T15108 = $signed(31'h3e44a5ee) * $signed(16'h1);
  assign twiddle4_2_39_real = T15114 + T15109;
  assign T15109 = {T15112, T15110};
  assign T15110 = $signed(T15111) / $signed(22'h100000);
  assign T15111 = $signed(29'hf2b650f) * $signed(16'h0);
  assign T15112 = T15113 ? 2'h3 : 2'h0;
  assign T15113 = T15110[6'h2c:6'h2c];
  assign T15114 = $signed(T15115) / $signed(22'h100000);
  assign T15115 = $signed(31'h3e2d1ea7) * $signed(16'h1);
  assign T15116 = T10817[1'h0:1'h0];
  assign T15117 = T10817[1'h1:1'h1];
  assign T15118 = T10817[2'h2:2'h2];
  assign T15119 = T15182 ? T15152 : T15120;
  assign T15120 = T15151 ? T15137 : T15121;
  assign T15121 = T15136 ? twiddle4_2_41_real : twiddle4_2_40_real;
  assign twiddle4_2_40_real = T15127 + T15122;
  assign T15122 = {T15125, T15123};
  assign T15123 = $signed(T15124) / $signed(22'h100000);
  assign T15124 = $signed(29'hf8cfcbd) * $signed(16'h0);
  assign T15125 = T15126 ? 2'h3 : 2'h0;
  assign T15126 = T15123[6'h2c:6'h2c];
  assign T15127 = $signed(T15128) / $signed(22'h100000);
  assign T15128 = $signed(31'h3e14fdf7) * $signed(16'h1);
  assign twiddle4_2_41_real = T15134 + T15129;
  assign T15129 = {T15132, T15130};
  assign T15130 = $signed(T15131) / $signed(22'h100000);
  assign T15131 = $signed(29'hfee6e0d) * $signed(16'h0);
  assign T15132 = T15133 ? 2'h3 : 2'h0;
  assign T15133 = T15130[6'h2c:6'h2c];
  assign T15134 = $signed(T15135) / $signed(22'h100000);
  assign T15135 = $signed(31'h3dfc4418) * $signed(16'h1);
  assign T15136 = T10817[1'h0:1'h0];
  assign T15137 = T15150 ? twiddle4_2_43_real : twiddle4_2_42_real;
  assign twiddle4_2_42_real = T15142 + T15138;
  assign T15138 = {T15141, T15139};
  assign T15139 = $signed(T15140) / $signed(22'h100000);
  assign T15140 = $signed(30'h104fb80e) * $signed(16'h0);
  assign T15141 = T15139[6'h2d:6'h2d];
  assign T15142 = $signed(T15143) / $signed(22'h100000);
  assign T15143 = $signed(31'h3de2f147) * $signed(16'h1);
  assign twiddle4_2_43_real = T15148 + T15144;
  assign T15144 = {T15147, T15145};
  assign T15145 = $signed(T15146) / $signed(22'h100000);
  assign T15146 = $signed(30'h10b0d9cf) * $signed(16'h0);
  assign T15147 = T15145[6'h2d:6'h2d];
  assign T15148 = $signed(T15149) / $signed(22'h100000);
  assign T15149 = $signed(31'h3dc905c4) * $signed(16'h1);
  assign T15150 = T10817[1'h0:1'h0];
  assign T15151 = T10817[1'h1:1'h1];
  assign T15152 = T15181 ? T15167 : T15153;
  assign T15153 = T15166 ? twiddle4_2_45_real : twiddle4_2_44_real;
  assign twiddle4_2_44_real = T15158 + T15154;
  assign T15154 = {T15157, T15155};
  assign T15155 = $signed(T15156) / $signed(22'h100000);
  assign T15156 = $signed(30'h1111d262) * $signed(16'h0);
  assign T15157 = T15155[6'h2d:6'h2d];
  assign T15158 = $signed(T15159) / $signed(22'h100000);
  assign T15159 = $signed(31'h3dae81ce) * $signed(16'h1);
  assign twiddle4_2_45_real = T15164 + T15160;
  assign T15160 = {T15163, T15161};
  assign T15161 = $signed(T15162) / $signed(22'h100000);
  assign T15162 = $signed(30'h1172a0d7) * $signed(16'h0);
  assign T15163 = T15161[6'h2d:6'h2d];
  assign T15164 = $signed(T15165) / $signed(22'h100000);
  assign T15165 = $signed(31'h3d9365a7) * $signed(16'h1);
  assign T15166 = T10817[1'h0:1'h0];
  assign T15167 = T15180 ? twiddle4_2_47_real : twiddle4_2_46_real;
  assign twiddle4_2_46_real = T15172 + T15168;
  assign T15168 = {T15171, T15169};
  assign T15169 = $signed(T15170) / $signed(22'h100000);
  assign T15170 = $signed(30'h11d3443f) * $signed(16'h0);
  assign T15171 = T15169[6'h2d:6'h2d];
  assign T15172 = $signed(T15173) / $signed(22'h100000);
  assign T15173 = $signed(31'h3d77b191) * $signed(16'h1);
  assign twiddle4_2_47_real = T15178 + T15174;
  assign T15174 = {T15177, T15175};
  assign T15175 = $signed(T15176) / $signed(22'h100000);
  assign T15176 = $signed(30'h1233bbab) * $signed(16'h0);
  assign T15177 = T15175[6'h2d:6'h2d];
  assign T15178 = $signed(T15179) / $signed(22'h100000);
  assign T15179 = $signed(31'h3d5b65d1) * $signed(16'h1);
  assign T15180 = T10817[1'h0:1'h0];
  assign T15181 = T10817[1'h1:1'h1];
  assign T15182 = T10817[2'h2:2'h2];
  assign T15183 = T10817[2'h3:2'h3];
  assign T15184 = T15309 ? T15247 : T15185;
  assign T15185 = T15246 ? T15216 : T15186;
  assign T15186 = T15215 ? T15201 : T15187;
  assign T15187 = T15200 ? twiddle4_2_49_real : twiddle4_2_48_real;
  assign twiddle4_2_48_real = T15192 + T15188;
  assign T15188 = {T15191, T15189};
  assign T15189 = $signed(T15190) / $signed(22'h100000);
  assign T15190 = $signed(30'h1294062e) * $signed(16'h0);
  assign T15191 = T15189[6'h2d:6'h2d];
  assign T15192 = $signed(T15193) / $signed(22'h100000);
  assign T15193 = $signed(31'h3d3e82ad) * $signed(16'h1);
  assign twiddle4_2_49_real = T15198 + T15194;
  assign T15194 = {T15197, T15195};
  assign T15195 = $signed(T15196) / $signed(22'h100000);
  assign T15196 = $signed(30'h12f422da) * $signed(16'h0);
  assign T15197 = T15195[6'h2d:6'h2d];
  assign T15198 = $signed(T15199) / $signed(22'h100000);
  assign T15199 = $signed(31'h3d21086c) * $signed(16'h1);
  assign T15200 = T10817[1'h0:1'h0];
  assign T15201 = T15214 ? twiddle4_2_51_real : twiddle4_2_50_real;
  assign twiddle4_2_50_real = T15206 + T15202;
  assign T15202 = {T15205, T15203};
  assign T15203 = $signed(T15204) / $signed(22'h100000);
  assign T15204 = $signed(30'h135410c2) * $signed(16'h0);
  assign T15205 = T15203[6'h2d:6'h2d];
  assign T15206 = $signed(T15207) / $signed(22'h100000);
  assign T15207 = $signed(31'h3d02f756) * $signed(16'h1);
  assign twiddle4_2_51_real = T15212 + T15208;
  assign T15208 = {T15211, T15209};
  assign T15209 = $signed(T15210) / $signed(22'h100000);
  assign T15210 = $signed(30'h13b3cefa) * $signed(16'h0);
  assign T15211 = T15209[6'h2d:6'h2d];
  assign T15212 = $signed(T15213) / $signed(22'h100000);
  assign T15213 = $signed(31'h3ce44fb6) * $signed(16'h1);
  assign T15214 = T10817[1'h0:1'h0];
  assign T15215 = T10817[1'h1:1'h1];
  assign T15216 = T15245 ? T15231 : T15217;
  assign T15217 = T15230 ? twiddle4_2_53_real : twiddle4_2_52_real;
  assign twiddle4_2_52_real = T15222 + T15218;
  assign T15218 = {T15221, T15219};
  assign T15219 = $signed(T15220) / $signed(22'h100000);
  assign T15220 = $signed(30'h14135c94) * $signed(16'h0);
  assign T15221 = T15219[6'h2d:6'h2d];
  assign T15222 = $signed(T15223) / $signed(22'h100000);
  assign T15223 = $signed(31'h3cc511d8) * $signed(16'h1);
  assign twiddle4_2_53_real = T15228 + T15224;
  assign T15224 = {T15227, T15225};
  assign T15225 = $signed(T15226) / $signed(22'h100000);
  assign T15226 = $signed(30'h1472b8a5) * $signed(16'h0);
  assign T15227 = T15225[6'h2d:6'h2d];
  assign T15228 = $signed(T15229) / $signed(22'h100000);
  assign T15229 = $signed(31'h3ca53e08) * $signed(16'h1);
  assign T15230 = T10817[1'h0:1'h0];
  assign T15231 = T15244 ? twiddle4_2_55_real : twiddle4_2_54_real;
  assign twiddle4_2_54_real = T15236 + T15232;
  assign T15232 = {T15235, T15233};
  assign T15233 = $signed(T15234) / $signed(22'h100000);
  assign T15234 = $signed(30'h14d1e242) * $signed(16'h0);
  assign T15235 = T15233[6'h2d:6'h2d];
  assign T15236 = $signed(T15237) / $signed(22'h100000);
  assign T15237 = $signed(31'h3c84d496) * $signed(16'h1);
  assign twiddle4_2_55_real = T15242 + T15238;
  assign T15238 = {T15241, T15239};
  assign T15239 = $signed(T15240) / $signed(22'h100000);
  assign T15240 = $signed(30'h1530d880) * $signed(16'h0);
  assign T15241 = T15239[6'h2d:6'h2d];
  assign T15242 = $signed(T15243) / $signed(22'h100000);
  assign T15243 = $signed(31'h3c63d5d0) * $signed(16'h1);
  assign T15244 = T10817[1'h0:1'h0];
  assign T15245 = T10817[1'h1:1'h1];
  assign T15246 = T10817[2'h2:2'h2];
  assign T15247 = T15308 ? T15278 : T15248;
  assign T15248 = T15277 ? T15263 : T15249;
  assign T15249 = T15262 ? twiddle4_2_57_real : twiddle4_2_56_real;
  assign twiddle4_2_56_real = T15254 + T15250;
  assign T15250 = {T15253, T15251};
  assign T15251 = $signed(T15252) / $signed(22'h100000);
  assign T15252 = $signed(30'h158f9a75) * $signed(16'h0);
  assign T15253 = T15251[6'h2d:6'h2d];
  assign T15254 = $signed(T15255) / $signed(22'h100000);
  assign T15255 = $signed(31'h3c424209) * $signed(16'h1);
  assign twiddle4_2_57_real = T15260 + T15256;
  assign T15256 = {T15259, T15257};
  assign T15257 = $signed(T15258) / $signed(22'h100000);
  assign T15258 = $signed(30'h15ee2737) * $signed(16'h0);
  assign T15259 = T15257[6'h2d:6'h2d];
  assign T15260 = $signed(T15261) / $signed(22'h100000);
  assign T15261 = $signed(31'h3c201994) * $signed(16'h1);
  assign T15262 = T10817[1'h0:1'h0];
  assign T15263 = T15276 ? twiddle4_2_59_real : twiddle4_2_58_real;
  assign twiddle4_2_58_real = T15268 + T15264;
  assign T15264 = {T15267, T15265};
  assign T15265 = $signed(T15266) / $signed(22'h100000);
  assign T15266 = $signed(30'h164c7ddd) * $signed(16'h0);
  assign T15267 = T15265[6'h2d:6'h2d];
  assign T15268 = $signed(T15269) / $signed(22'h100000);
  assign T15269 = $signed(31'h3bfd5cc4) * $signed(16'h1);
  assign twiddle4_2_59_real = T15274 + T15270;
  assign T15270 = {T15273, T15271};
  assign T15271 = $signed(T15272) / $signed(22'h100000);
  assign T15272 = $signed(30'h16aa9d7d) * $signed(16'h0);
  assign T15273 = T15271[6'h2d:6'h2d];
  assign T15274 = $signed(T15275) / $signed(22'h100000);
  assign T15275 = $signed(31'h3bda0bef) * $signed(16'h1);
  assign T15276 = T10817[1'h0:1'h0];
  assign T15277 = T10817[1'h1:1'h1];
  assign T15278 = T15307 ? T15293 : T15279;
  assign T15279 = T15292 ? twiddle4_2_61_real : twiddle4_2_60_real;
  assign twiddle4_2_60_real = T15284 + T15280;
  assign T15280 = {T15283, T15281};
  assign T15281 = $signed(T15282) / $signed(22'h100000);
  assign T15282 = $signed(30'h17088530) * $signed(16'h0);
  assign T15283 = T15281[6'h2d:6'h2d];
  assign T15284 = $signed(T15285) / $signed(22'h100000);
  assign T15285 = $signed(31'h3bb6276d) * $signed(16'h1);
  assign twiddle4_2_61_real = T15290 + T15286;
  assign T15286 = {T15289, T15287};
  assign T15287 = $signed(T15288) / $signed(22'h100000);
  assign T15288 = $signed(30'h1766340f) * $signed(16'h0);
  assign T15289 = T15287[6'h2d:6'h2d];
  assign T15290 = $signed(T15291) / $signed(22'h100000);
  assign T15291 = $signed(31'h3b91af96) * $signed(16'h1);
  assign T15292 = T10817[1'h0:1'h0];
  assign T15293 = T15306 ? twiddle4_2_63_real : twiddle4_2_62_real;
  assign twiddle4_2_62_real = T15298 + T15294;
  assign T15294 = {T15297, T15295};
  assign T15295 = $signed(T15296) / $signed(22'h100000);
  assign T15296 = $signed(30'h17c3a931) * $signed(16'h0);
  assign T15297 = T15295[6'h2d:6'h2d];
  assign T15298 = $signed(T15299) / $signed(22'h100000);
  assign T15299 = $signed(31'h3b6ca4c4) * $signed(16'h1);
  assign twiddle4_2_63_real = T15304 + T15300;
  assign T15300 = {T15303, T15301};
  assign T15301 = $signed(T15302) / $signed(22'h100000);
  assign T15302 = $signed(30'h1820e3b0) * $signed(16'h0);
  assign T15303 = T15301[6'h2d:6'h2d];
  assign T15304 = $signed(T15305) / $signed(22'h100000);
  assign T15305 = $signed(31'h3b470752) * $signed(16'h1);
  assign T15306 = T10817[1'h0:1'h0];
  assign T15307 = T10817[1'h1:1'h1];
  assign T15308 = T10817[2'h2:2'h2];
  assign T15309 = T10817[2'h3:2'h3];
  assign T15310 = T10817[3'h4:3'h4];
  assign T15311 = T15047[6'h2e:6'h2e];
  assign T15312 = T10817[3'h5:3'h5];
  assign T15313 = {T15740, T15314};
  assign T15314 = T15739 ? T15549 : T15315;
  assign T15315 = T15548 ? T15442 : T15316;
  assign T15316 = T15441 ? T15379 : T15317;
  assign T15317 = T15378 ? T15348 : T15318;
  assign T15318 = T15347 ? T15333 : T15319;
  assign T15319 = T15332 ? twiddle4_2_65_real : twiddle4_2_64_real;
  assign twiddle4_2_64_real = T15324 + T15320;
  assign T15320 = {T15323, T15321};
  assign T15321 = $signed(T15322) / $signed(22'h100000);
  assign T15322 = $signed(30'h187de2a6) * $signed(16'h0);
  assign T15323 = T15321[6'h2d:6'h2d];
  assign T15324 = $signed(T15325) / $signed(22'h100000);
  assign T15325 = $signed(31'h3b20d79e) * $signed(16'h1);
  assign twiddle4_2_65_real = T15330 + T15326;
  assign T15326 = {T15329, T15327};
  assign T15327 = $signed(T15328) / $signed(22'h100000);
  assign T15328 = $signed(30'h18daa52e) * $signed(16'h0);
  assign T15329 = T15327[6'h2d:6'h2d];
  assign T15330 = $signed(T15331) / $signed(22'h100000);
  assign T15331 = $signed(31'h3afa1605) * $signed(16'h1);
  assign T15332 = T10817[1'h0:1'h0];
  assign T15333 = T15346 ? twiddle4_2_67_real : twiddle4_2_66_real;
  assign twiddle4_2_66_real = T15338 + T15334;
  assign T15334 = {T15337, T15335};
  assign T15335 = $signed(T15336) / $signed(22'h100000);
  assign T15336 = $signed(30'h19372a63) * $signed(16'h0);
  assign T15337 = T15335[6'h2d:6'h2d];
  assign T15338 = $signed(T15339) / $signed(22'h100000);
  assign T15339 = $signed(31'h3ad2c2e7) * $signed(16'h1);
  assign twiddle4_2_67_real = T15344 + T15340;
  assign T15340 = {T15343, T15341};
  assign T15341 = $signed(T15342) / $signed(22'h100000);
  assign T15342 = $signed(30'h19937161) * $signed(16'h0);
  assign T15343 = T15341[6'h2d:6'h2d];
  assign T15344 = $signed(T15345) / $signed(22'h100000);
  assign T15345 = $signed(31'h3aaadea5) * $signed(16'h1);
  assign T15346 = T10817[1'h0:1'h0];
  assign T15347 = T10817[1'h1:1'h1];
  assign T15348 = T15377 ? T15363 : T15349;
  assign T15349 = T15362 ? twiddle4_2_69_real : twiddle4_2_68_real;
  assign twiddle4_2_68_real = T15354 + T15350;
  assign T15350 = {T15353, T15351};
  assign T15351 = $signed(T15352) / $signed(22'h100000);
  assign T15352 = $signed(30'h19ef7943) * $signed(16'h0);
  assign T15353 = T15351[6'h2d:6'h2d];
  assign T15354 = $signed(T15355) / $signed(22'h100000);
  assign T15355 = $signed(31'h3a8269a2) * $signed(16'h1);
  assign twiddle4_2_69_real = T15360 + T15356;
  assign T15356 = {T15359, T15357};
  assign T15357 = $signed(T15358) / $signed(22'h100000);
  assign T15358 = $signed(30'h1a4b4127) * $signed(16'h0);
  assign T15359 = T15357[6'h2d:6'h2d];
  assign T15360 = $signed(T15361) / $signed(22'h100000);
  assign T15361 = $signed(31'h3a596441) * $signed(16'h1);
  assign T15362 = T10817[1'h0:1'h0];
  assign T15363 = T15376 ? twiddle4_2_71_real : twiddle4_2_70_real;
  assign twiddle4_2_70_real = T15368 + T15364;
  assign T15364 = {T15367, T15365};
  assign T15365 = $signed(T15366) / $signed(22'h100000);
  assign T15366 = $signed(30'h1aa6c82b) * $signed(16'h0);
  assign T15367 = T15365[6'h2d:6'h2d];
  assign T15368 = $signed(T15369) / $signed(22'h100000);
  assign T15369 = $signed(31'h3a2fcee8) * $signed(16'h1);
  assign twiddle4_2_71_real = T15374 + T15370;
  assign T15370 = {T15373, T15371};
  assign T15371 = $signed(T15372) / $signed(22'h100000);
  assign T15372 = $signed(30'h1b020d6c) * $signed(16'h0);
  assign T15373 = T15371[6'h2d:6'h2d];
  assign T15374 = $signed(T15375) / $signed(22'h100000);
  assign T15375 = $signed(31'h3a05a9fd) * $signed(16'h1);
  assign T15376 = T10817[1'h0:1'h0];
  assign T15377 = T10817[1'h1:1'h1];
  assign T15378 = T10817[2'h2:2'h2];
  assign T15379 = T15440 ? T15410 : T15380;
  assign T15380 = T15409 ? T15395 : T15381;
  assign T15381 = T15394 ? twiddle4_2_73_real : twiddle4_2_72_real;
  assign twiddle4_2_72_real = T15386 + T15382;
  assign T15382 = {T15385, T15383};
  assign T15383 = $signed(T15384) / $signed(22'h100000);
  assign T15384 = $signed(30'h1b5d1009) * $signed(16'h0);
  assign T15385 = T15383[6'h2d:6'h2d];
  assign T15386 = $signed(T15387) / $signed(22'h100000);
  assign T15387 = $signed(31'h39daf5e8) * $signed(16'h1);
  assign twiddle4_2_73_real = T15392 + T15388;
  assign T15388 = {T15391, T15389};
  assign T15389 = $signed(T15390) / $signed(22'h100000);
  assign T15390 = $signed(30'h1bb7cf23) * $signed(16'h0);
  assign T15391 = T15389[6'h2d:6'h2d];
  assign T15392 = $signed(T15393) / $signed(22'h100000);
  assign T15393 = $signed(31'h39afb313) * $signed(16'h1);
  assign T15394 = T10817[1'h0:1'h0];
  assign T15395 = T15408 ? twiddle4_2_75_real : twiddle4_2_74_real;
  assign twiddle4_2_74_real = T15400 + T15396;
  assign T15396 = {T15399, T15397};
  assign T15397 = $signed(T15398) / $signed(22'h100000);
  assign T15398 = $signed(30'h1c1249d8) * $signed(16'h0);
  assign T15399 = T15397[6'h2d:6'h2d];
  assign T15400 = $signed(T15401) / $signed(22'h100000);
  assign T15401 = $signed(31'h3983e1e7) * $signed(16'h1);
  assign twiddle4_2_75_real = T15406 + T15402;
  assign T15402 = {T15405, T15403};
  assign T15403 = $signed(T15404) / $signed(22'h100000);
  assign T15404 = $signed(30'h1c6c7f49) * $signed(16'h0);
  assign T15405 = T15403[6'h2d:6'h2d];
  assign T15406 = $signed(T15407) / $signed(22'h100000);
  assign T15407 = $signed(31'h395782d3) * $signed(16'h1);
  assign T15408 = T10817[1'h0:1'h0];
  assign T15409 = T10817[1'h1:1'h1];
  assign T15410 = T15439 ? T15425 : T15411;
  assign T15411 = T15424 ? twiddle4_2_77_real : twiddle4_2_76_real;
  assign twiddle4_2_76_real = T15416 + T15412;
  assign T15412 = {T15415, T15413};
  assign T15413 = $signed(T15414) / $signed(22'h100000);
  assign T15414 = $signed(30'h1cc66e99) * $signed(16'h0);
  assign T15415 = T15413[6'h2d:6'h2d];
  assign T15416 = $signed(T15417) / $signed(22'h100000);
  assign T15417 = $signed(31'h392a9642) * $signed(16'h1);
  assign twiddle4_2_77_real = T15422 + T15418;
  assign T15418 = {T15421, T15419};
  assign T15419 = $signed(T15420) / $signed(22'h100000);
  assign T15420 = $signed(30'h1d2016e8) * $signed(16'h0);
  assign T15421 = T15419[6'h2d:6'h2d];
  assign T15422 = $signed(T15423) / $signed(22'h100000);
  assign T15423 = $signed(31'h38fd1ca4) * $signed(16'h1);
  assign T15424 = T10817[1'h0:1'h0];
  assign T15425 = T15438 ? twiddle4_2_79_real : twiddle4_2_78_real;
  assign twiddle4_2_78_real = T15430 + T15426;
  assign T15426 = {T15429, T15427};
  assign T15427 = $signed(T15428) / $signed(22'h100000);
  assign T15428 = $signed(30'h1d79775b) * $signed(16'h0);
  assign T15429 = T15427[6'h2d:6'h2d];
  assign T15430 = $signed(T15431) / $signed(22'h100000);
  assign T15431 = $signed(31'h38cf1669) * $signed(16'h1);
  assign twiddle4_2_79_real = T15436 + T15432;
  assign T15432 = {T15435, T15433};
  assign T15433 = $signed(T15434) / $signed(22'h100000);
  assign T15434 = $signed(30'h1dd28f14) * $signed(16'h0);
  assign T15435 = T15433[6'h2d:6'h2d];
  assign T15436 = $signed(T15437) / $signed(22'h100000);
  assign T15437 = $signed(31'h38a08402) * $signed(16'h1);
  assign T15438 = T10817[1'h0:1'h0];
  assign T15439 = T10817[1'h1:1'h1];
  assign T15440 = T10817[2'h2:2'h2];
  assign T15441 = T10817[2'h3:2'h3];
  assign T15442 = T15547 ? T15501 : T15443;
  assign T15443 = T15500 ? T15474 : T15444;
  assign T15444 = T15473 ? T15459 : T15445;
  assign T15445 = T15458 ? twiddle4_2_81_real : twiddle4_2_80_real;
  assign twiddle4_2_80_real = T15450 + T15446;
  assign T15446 = {T15449, T15447};
  assign T15447 = $signed(T15448) / $signed(22'h100000);
  assign T15448 = $signed(30'h1e2b5d38) * $signed(16'h0);
  assign T15449 = T15447[6'h2d:6'h2d];
  assign T15450 = $signed(T15451) / $signed(22'h100000);
  assign T15451 = $signed(31'h387165e3) * $signed(16'h1);
  assign twiddle4_2_81_real = T15456 + T15452;
  assign T15452 = {T15455, T15453};
  assign T15453 = $signed(T15454) / $signed(22'h100000);
  assign T15454 = $signed(30'h1e83e0ea) * $signed(16'h0);
  assign T15455 = T15453[6'h2d:6'h2d];
  assign T15456 = $signed(T15457) / $signed(22'h100000);
  assign T15457 = $signed(31'h3841bc7f) * $signed(16'h1);
  assign T15458 = T10817[1'h0:1'h0];
  assign T15459 = T15472 ? twiddle4_2_83_real : twiddle4_2_82_real;
  assign twiddle4_2_82_real = T15464 + T15460;
  assign T15460 = {T15463, T15461};
  assign T15461 = $signed(T15462) / $signed(22'h100000);
  assign T15462 = $signed(30'h1edc1952) * $signed(16'h0);
  assign T15463 = T15461[6'h2d:6'h2d];
  assign T15464 = $signed(T15465) / $signed(22'h100000);
  assign T15465 = $signed(31'h3811884c) * $signed(16'h1);
  assign twiddle4_2_83_real = T15470 + T15466;
  assign T15466 = {T15469, T15467};
  assign T15467 = $signed(T15468) / $signed(22'h100000);
  assign T15468 = $signed(30'h1f340596) * $signed(16'h0);
  assign T15469 = T15467[6'h2d:6'h2d];
  assign T15470 = $signed(T15471) / $signed(22'h100000);
  assign T15471 = $signed(31'h37e0c9c2) * $signed(16'h1);
  assign T15472 = T10817[1'h0:1'h0];
  assign T15473 = T10817[1'h1:1'h1];
  assign T15474 = T15499 ? T15489 : T15475;
  assign T15475 = T15488 ? twiddle4_2_85_real : twiddle4_2_84_real;
  assign twiddle4_2_84_real = T15480 + T15476;
  assign T15476 = {T15479, T15477};
  assign T15477 = $signed(T15478) / $signed(22'h100000);
  assign T15478 = $signed(30'h1f8ba4db) * $signed(16'h0);
  assign T15479 = T15477[6'h2d:6'h2d];
  assign T15480 = $signed(T15481) / $signed(22'h100000);
  assign T15481 = $signed(31'h37af8158) * $signed(16'h1);
  assign twiddle4_2_85_real = T15486 + T15482;
  assign T15482 = {T15485, T15483};
  assign T15483 = $signed(T15484) / $signed(22'h100000);
  assign T15484 = $signed(30'h1fe2f64b) * $signed(16'h0);
  assign T15485 = T15483[6'h2d:6'h2d];
  assign T15486 = $signed(T15487) / $signed(22'h100000);
  assign T15487 = $signed(31'h377daf89) * $signed(16'h1);
  assign T15488 = T10817[1'h0:1'h0];
  assign T15489 = T15498 ? twiddle4_2_87_real : twiddle4_2_86_real;
  assign twiddle4_2_86_real = T15492 + T15490;
  assign T15490 = $signed(T15491) / $signed(22'h100000);
  assign T15491 = $signed(31'h2039f90e) * $signed(16'h0);
  assign T15492 = $signed(T15493) / $signed(22'h100000);
  assign T15493 = $signed(31'h374b54ce) * $signed(16'h1);
  assign twiddle4_2_87_real = T15496 + T15494;
  assign T15494 = $signed(T15495) / $signed(22'h100000);
  assign T15495 = $signed(31'h2090ac4d) * $signed(16'h0);
  assign T15496 = $signed(T15497) / $signed(22'h100000);
  assign T15497 = $signed(31'h371871a4) * $signed(16'h1);
  assign T15498 = T10817[1'h0:1'h0];
  assign T15499 = T10817[1'h1:1'h1];
  assign T15500 = T10817[2'h2:2'h2];
  assign T15501 = T15546 ? T15524 : T15502;
  assign T15502 = T15523 ? T15513 : T15503;
  assign T15503 = T15512 ? twiddle4_2_89_real : twiddle4_2_88_real;
  assign twiddle4_2_88_real = T15506 + T15504;
  assign T15504 = $signed(T15505) / $signed(22'h100000);
  assign T15505 = $signed(31'h20e70f32) * $signed(16'h0);
  assign T15506 = $signed(T15507) / $signed(22'h100000);
  assign T15507 = $signed(31'h36e5068a) * $signed(16'h1);
  assign twiddle4_2_89_real = T15510 + T15508;
  assign T15508 = $signed(T15509) / $signed(22'h100000);
  assign T15509 = $signed(31'h213d20e8) * $signed(16'h0);
  assign T15510 = $signed(T15511) / $signed(22'h100000);
  assign T15511 = $signed(31'h36b113fd) * $signed(16'h1);
  assign T15512 = T10817[1'h0:1'h0];
  assign T15513 = T15522 ? twiddle4_2_91_real : twiddle4_2_90_real;
  assign twiddle4_2_90_real = T15516 + T15514;
  assign T15514 = $signed(T15515) / $signed(22'h100000);
  assign T15515 = $signed(31'h2192e09a) * $signed(16'h0);
  assign T15516 = $signed(T15517) / $signed(22'h100000);
  assign T15517 = $signed(31'h367c9a7d) * $signed(16'h1);
  assign twiddle4_2_91_real = T15520 + T15518;
  assign T15518 = $signed(T15519) / $signed(22'h100000);
  assign T15519 = $signed(31'h21e84d76) * $signed(16'h0);
  assign T15520 = $signed(T15521) / $signed(22'h100000);
  assign T15521 = $signed(31'h36479a8e) * $signed(16'h1);
  assign T15522 = T10817[1'h0:1'h0];
  assign T15523 = T10817[1'h1:1'h1];
  assign T15524 = T15545 ? T15535 : T15525;
  assign T15525 = T15534 ? twiddle4_2_93_real : twiddle4_2_92_real;
  assign twiddle4_2_92_real = T15528 + T15526;
  assign T15526 = $signed(T15527) / $signed(22'h100000);
  assign T15527 = $signed(31'h223d66a8) * $signed(16'h0);
  assign T15528 = $signed(T15529) / $signed(22'h100000);
  assign T15529 = $signed(31'h361214b0) * $signed(16'h1);
  assign twiddle4_2_93_real = T15532 + T15530;
  assign T15530 = $signed(T15531) / $signed(22'h100000);
  assign T15531 = $signed(31'h22922b5e) * $signed(16'h0);
  assign T15532 = $signed(T15533) / $signed(22'h100000);
  assign T15533 = $signed(31'h35dc0968) * $signed(16'h1);
  assign T15534 = T10817[1'h0:1'h0];
  assign T15535 = T15544 ? twiddle4_2_95_real : twiddle4_2_94_real;
  assign twiddle4_2_94_real = T15538 + T15536;
  assign T15536 = $signed(T15537) / $signed(22'h100000);
  assign T15537 = $signed(31'h22e69ac7) * $signed(16'h0);
  assign T15538 = $signed(T15539) / $signed(22'h100000);
  assign T15539 = $signed(31'h35a5793c) * $signed(16'h1);
  assign twiddle4_2_95_real = T15542 + T15540;
  assign T15540 = $signed(T15541) / $signed(22'h100000);
  assign T15541 = $signed(31'h233ab413) * $signed(16'h0);
  assign T15542 = $signed(T15543) / $signed(22'h100000);
  assign T15543 = $signed(31'h356e64b2) * $signed(16'h1);
  assign T15544 = T10817[1'h0:1'h0];
  assign T15545 = T10817[1'h1:1'h1];
  assign T15546 = T10817[2'h2:2'h2];
  assign T15547 = T10817[2'h3:2'h3];
  assign T15548 = T10817[3'h4:3'h4];
  assign T15549 = T15738 ? T15644 : T15550;
  assign T15550 = T15643 ? T15597 : T15551;
  assign T15551 = T15596 ? T15574 : T15552;
  assign T15552 = T15573 ? T15563 : T15553;
  assign T15553 = T15562 ? twiddle4_2_97_real : twiddle4_2_96_real;
  assign twiddle4_2_96_real = T15556 + T15554;
  assign T15554 = $signed(T15555) / $signed(22'h100000);
  assign T15555 = $signed(31'h238e7673) * $signed(16'h0);
  assign T15556 = $signed(T15557) / $signed(22'h100000);
  assign T15557 = $signed(31'h3536cc52) * $signed(16'h1);
  assign twiddle4_2_97_real = T15560 + T15558;
  assign T15558 = $signed(T15559) / $signed(22'h100000);
  assign T15559 = $signed(31'h23e1e117) * $signed(16'h0);
  assign T15560 = $signed(T15561) / $signed(22'h100000);
  assign T15561 = $signed(31'h34feb0a5) * $signed(16'h1);
  assign T15562 = T10817[1'h0:1'h0];
  assign T15563 = T15572 ? twiddle4_2_99_real : twiddle4_2_98_real;
  assign twiddle4_2_98_real = T15566 + T15564;
  assign T15564 = $signed(T15565) / $signed(22'h100000);
  assign T15565 = $signed(31'h2434f332) * $signed(16'h0);
  assign T15566 = $signed(T15567) / $signed(22'h100000);
  assign T15567 = $signed(31'h34c61236) * $signed(16'h1);
  assign twiddle4_2_99_real = T15570 + T15568;
  assign T15568 = $signed(T15569) / $signed(22'h100000);
  assign T15569 = $signed(31'h2487abf7) * $signed(16'h0);
  assign T15570 = $signed(T15571) / $signed(22'h100000);
  assign T15571 = $signed(31'h348cf190) * $signed(16'h1);
  assign T15572 = T10817[1'h0:1'h0];
  assign T15573 = T10817[1'h1:1'h1];
  assign T15574 = T15595 ? T15585 : T15575;
  assign T15575 = T15584 ? twiddle4_2_101_real : twiddle4_2_100_real;
  assign twiddle4_2_100_real = T15578 + T15576;
  assign T15576 = $signed(T15577) / $signed(22'h100000);
  assign T15577 = $signed(31'h24da0a99) * $signed(16'h0);
  assign T15578 = $signed(T15579) / $signed(22'h100000);
  assign T15579 = $signed(31'h34534f40) * $signed(16'h1);
  assign twiddle4_2_101_real = T15582 + T15580;
  assign T15580 = $signed(T15581) / $signed(22'h100000);
  assign T15581 = $signed(31'h252c0e4e) * $signed(16'h0);
  assign T15582 = $signed(T15583) / $signed(22'h100000);
  assign T15583 = $signed(31'h34192bd5) * $signed(16'h1);
  assign T15584 = T10817[1'h0:1'h0];
  assign T15585 = T15594 ? twiddle4_2_103_real : twiddle4_2_102_real;
  assign twiddle4_2_102_real = T15588 + T15586;
  assign T15586 = $signed(T15587) / $signed(22'h100000);
  assign T15587 = $signed(31'h257db64b) * $signed(16'h0);
  assign T15588 = $signed(T15589) / $signed(22'h100000);
  assign T15589 = $signed(31'h33de87de) * $signed(16'h1);
  assign twiddle4_2_103_real = T15592 + T15590;
  assign T15590 = $signed(T15591) / $signed(22'h100000);
  assign T15591 = $signed(31'h25cf01c7) * $signed(16'h0);
  assign T15592 = $signed(T15593) / $signed(22'h100000);
  assign T15593 = $signed(31'h33a363eb) * $signed(16'h1);
  assign T15594 = T10817[1'h0:1'h0];
  assign T15595 = T10817[1'h1:1'h1];
  assign T15596 = T10817[2'h2:2'h2];
  assign T15597 = T15642 ? T15620 : T15598;
  assign T15598 = T15619 ? T15609 : T15599;
  assign T15599 = T15608 ? twiddle4_2_105_real : twiddle4_2_104_real;
  assign twiddle4_2_104_real = T15602 + T15600;
  assign T15600 = $signed(T15601) / $signed(22'h100000);
  assign T15601 = $signed(31'h261feff9) * $signed(16'h0);
  assign T15602 = $signed(T15603) / $signed(22'h100000);
  assign T15603 = $signed(31'h3367c08f) * $signed(16'h1);
  assign twiddle4_2_105_real = T15606 + T15604;
  assign T15604 = $signed(T15605) / $signed(22'h100000);
  assign T15605 = $signed(31'h2670801a) * $signed(16'h0);
  assign T15606 = $signed(T15607) / $signed(22'h100000);
  assign T15607 = $signed(31'h332b9e5d) * $signed(16'h1);
  assign T15608 = T10817[1'h0:1'h0];
  assign T15609 = T15618 ? twiddle4_2_107_real : twiddle4_2_106_real;
  assign twiddle4_2_106_real = T15612 + T15610;
  assign T15610 = $signed(T15611) / $signed(22'h100000);
  assign T15611 = $signed(31'h26c0b162) * $signed(16'h0);
  assign T15612 = $signed(T15613) / $signed(22'h100000);
  assign T15613 = $signed(31'h32eefde9) * $signed(16'h1);
  assign twiddle4_2_107_real = T15616 + T15614;
  assign T15614 = $signed(T15615) / $signed(22'h100000);
  assign T15615 = $signed(31'h2710830b) * $signed(16'h0);
  assign T15616 = $signed(T15617) / $signed(22'h100000);
  assign T15617 = $signed(31'h32b1dfc9) * $signed(16'h1);
  assign T15618 = T10817[1'h0:1'h0];
  assign T15619 = T10817[1'h1:1'h1];
  assign T15620 = T15641 ? T15631 : T15621;
  assign T15621 = T15630 ? twiddle4_2_109_real : twiddle4_2_108_real;
  assign twiddle4_2_108_real = T15624 + T15622;
  assign T15622 = $signed(T15623) / $signed(22'h100000);
  assign T15623 = $signed(31'h275ff452) * $signed(16'h0);
  assign T15624 = $signed(T15625) / $signed(22'h100000);
  assign T15625 = $signed(31'h32744493) * $signed(16'h1);
  assign twiddle4_2_109_real = T15628 + T15626;
  assign T15626 = $signed(T15627) / $signed(22'h100000);
  assign T15627 = $signed(31'h27af0471) * $signed(16'h0);
  assign T15628 = $signed(T15629) / $signed(22'h100000);
  assign T15629 = $signed(31'h32362cdf) * $signed(16'h1);
  assign T15630 = T10817[1'h0:1'h0];
  assign T15631 = T15640 ? twiddle4_2_111_real : twiddle4_2_110_real;
  assign twiddle4_2_110_real = T15634 + T15632;
  assign T15632 = $signed(T15633) / $signed(22'h100000);
  assign T15633 = $signed(31'h27fdb2a6) * $signed(16'h0);
  assign T15634 = $signed(T15635) / $signed(22'h100000);
  assign T15635 = $signed(31'h31f79947) * $signed(16'h1);
  assign twiddle4_2_111_real = T15638 + T15636;
  assign T15636 = $signed(T15637) / $signed(22'h100000);
  assign T15637 = $signed(31'h284bfe2f) * $signed(16'h0);
  assign T15638 = $signed(T15639) / $signed(22'h100000);
  assign T15639 = $signed(31'h31b88a66) * $signed(16'h1);
  assign T15640 = T10817[1'h0:1'h0];
  assign T15641 = T10817[1'h1:1'h1];
  assign T15642 = T10817[2'h2:2'h2];
  assign T15643 = T10817[2'h3:2'h3];
  assign T15644 = T15737 ? T15691 : T15645;
  assign T15645 = T15690 ? T15668 : T15646;
  assign T15646 = T15667 ? T15657 : T15647;
  assign T15647 = T15656 ? twiddle4_2_113_real : twiddle4_2_112_real;
  assign twiddle4_2_112_real = T15650 + T15648;
  assign T15648 = $signed(T15649) / $signed(22'h100000);
  assign T15649 = $signed(31'h2899e64a) * $signed(16'h0);
  assign T15650 = $signed(T15651) / $signed(22'h100000);
  assign T15651 = $signed(31'h317900d6) * $signed(16'h1);
  assign twiddle4_2_113_real = T15654 + T15652;
  assign T15652 = $signed(T15653) / $signed(22'h100000);
  assign T15653 = $signed(31'h28e76a37) * $signed(16'h0);
  assign T15654 = $signed(T15655) / $signed(22'h100000);
  assign T15655 = $signed(31'h3138fd34) * $signed(16'h1);
  assign T15656 = T10817[1'h0:1'h0];
  assign T15657 = T15666 ? twiddle4_2_115_real : twiddle4_2_114_real;
  assign twiddle4_2_114_real = T15660 + T15658;
  assign T15658 = $signed(T15659) / $signed(22'h100000);
  assign T15659 = $signed(31'h29348937) * $signed(16'h0);
  assign T15660 = $signed(T15661) / $signed(22'h100000);
  assign T15661 = $signed(31'h30f8801f) * $signed(16'h1);
  assign twiddle4_2_115_real = T15664 + T15662;
  assign T15662 = $signed(T15663) / $signed(22'h100000);
  assign T15663 = $signed(31'h2981428b) * $signed(16'h0);
  assign T15664 = $signed(T15665) / $signed(22'h100000);
  assign T15665 = $signed(31'h30b78a35) * $signed(16'h1);
  assign T15666 = T10817[1'h0:1'h0];
  assign T15667 = T10817[1'h1:1'h1];
  assign T15668 = T15689 ? T15679 : T15669;
  assign T15669 = T15678 ? twiddle4_2_117_real : twiddle4_2_116_real;
  assign twiddle4_2_116_real = T15672 + T15670;
  assign T15670 = $signed(T15671) / $signed(22'h100000);
  assign T15671 = $signed(31'h29cd9577) * $signed(16'h0);
  assign T15672 = $signed(T15673) / $signed(22'h100000);
  assign T15673 = $signed(31'h30761c17) * $signed(16'h1);
  assign twiddle4_2_117_real = T15676 + T15674;
  assign T15674 = $signed(T15675) / $signed(22'h100000);
  assign T15675 = $signed(31'h2a19813e) * $signed(16'h0);
  assign T15676 = $signed(T15677) / $signed(22'h100000);
  assign T15677 = $signed(31'h30343667) * $signed(16'h1);
  assign T15678 = T10817[1'h0:1'h0];
  assign T15679 = T15688 ? twiddle4_2_119_real : twiddle4_2_118_real;
  assign twiddle4_2_118_real = T15682 + T15680;
  assign T15680 = $signed(T15681) / $signed(22'h100000);
  assign T15681 = $signed(31'h2a650525) * $signed(16'h0);
  assign T15682 = $signed(T15683) / $signed(22'h100000);
  assign T15683 = $signed(31'h2ff1d9c6) * $signed(16'h1);
  assign twiddle4_2_119_real = T15686 + T15684;
  assign T15684 = $signed(T15685) / $signed(22'h100000);
  assign T15685 = $signed(31'h2ab02071) * $signed(16'h0);
  assign T15686 = $signed(T15687) / $signed(22'h100000);
  assign T15687 = $signed(31'h2faf06d9) * $signed(16'h1);
  assign T15688 = T10817[1'h0:1'h0];
  assign T15689 = T10817[1'h1:1'h1];
  assign T15690 = T10817[2'h2:2'h2];
  assign T15691 = T15736 ? T15714 : T15692;
  assign T15692 = T15713 ? T15703 : T15693;
  assign T15693 = T15702 ? twiddle4_2_121_real : twiddle4_2_120_real;
  assign twiddle4_2_120_real = T15696 + T15694;
  assign T15694 = $signed(T15695) / $signed(22'h100000);
  assign T15695 = $signed(31'h2afad269) * $signed(16'h0);
  assign T15696 = $signed(T15697) / $signed(22'h100000);
  assign T15697 = $signed(31'h2f6bbe44) * $signed(16'h1);
  assign twiddle4_2_121_real = T15700 + T15698;
  assign T15698 = $signed(T15699) / $signed(22'h100000);
  assign T15699 = $signed(31'h2b451a54) * $signed(16'h0);
  assign T15700 = $signed(T15701) / $signed(22'h100000);
  assign T15701 = $signed(31'h2f2800ae) * $signed(16'h1);
  assign T15702 = T10817[1'h0:1'h0];
  assign T15703 = T15712 ? twiddle4_2_123_real : twiddle4_2_122_real;
  assign twiddle4_2_122_real = T15706 + T15704;
  assign T15704 = $signed(T15705) / $signed(22'h100000);
  assign T15705 = $signed(31'h2b8ef77c) * $signed(16'h0);
  assign T15706 = $signed(T15707) / $signed(22'h100000);
  assign T15707 = $signed(31'h2ee3cebe) * $signed(16'h1);
  assign twiddle4_2_123_real = T15710 + T15708;
  assign T15708 = $signed(T15709) / $signed(22'h100000);
  assign T15709 = $signed(31'h2bd8692b) * $signed(16'h0);
  assign T15710 = $signed(T15711) / $signed(22'h100000);
  assign T15711 = $signed(31'h2e9f291b) * $signed(16'h1);
  assign T15712 = T10817[1'h0:1'h0];
  assign T15713 = T10817[1'h1:1'h1];
  assign T15714 = T15735 ? T15725 : T15715;
  assign T15715 = T15724 ? twiddle4_2_125_real : twiddle4_2_124_real;
  assign twiddle4_2_124_real = T15718 + T15716;
  assign T15716 = $signed(T15717) / $signed(22'h100000);
  assign T15717 = $signed(31'h2c216eaa) * $signed(16'h0);
  assign T15718 = $signed(T15719) / $signed(22'h100000);
  assign T15719 = $signed(31'h2e5a106f) * $signed(16'h1);
  assign twiddle4_2_125_real = T15722 + T15720;
  assign T15720 = $signed(T15721) / $signed(22'h100000);
  assign T15721 = $signed(31'h2c6a0746) * $signed(16'h0);
  assign T15722 = $signed(T15723) / $signed(22'h100000);
  assign T15723 = $signed(31'h2e148566) * $signed(16'h1);
  assign T15724 = T10817[1'h0:1'h0];
  assign T15725 = T15734 ? twiddle4_2_127_real : twiddle4_2_126_real;
  assign twiddle4_2_126_real = T15728 + T15726;
  assign T15726 = $signed(T15727) / $signed(22'h100000);
  assign T15727 = $signed(31'h2cb2324b) * $signed(16'h0);
  assign T15728 = $signed(T15729) / $signed(22'h100000);
  assign T15729 = $signed(31'h2dce88a9) * $signed(16'h1);
  assign twiddle4_2_127_real = T15732 + T15730;
  assign T15730 = $signed(T15731) / $signed(22'h100000);
  assign T15731 = $signed(31'h2cf9ef09) * $signed(16'h0);
  assign T15732 = $signed(T15733) / $signed(22'h100000);
  assign T15733 = $signed(31'h2d881ae7) * $signed(16'h1);
  assign T15734 = T10817[1'h0:1'h0];
  assign T15735 = T10817[1'h1:1'h1];
  assign T15736 = T10817[2'h2:2'h2];
  assign T15737 = T10817[2'h3:2'h3];
  assign T15738 = T10817[3'h4:3'h4];
  assign T15739 = T10817[3'h5:3'h5];
  assign T15740 = T15314[6'h2e:6'h2e];
  assign T15741 = T10817[3'h6:3'h6];
  assign T15742 = {T16720, T15743};
  assign T15743 = T16719 ? T16168 : T15744;
  assign T15744 = T16167 ? T15935 : T15745;
  assign T15745 = T15934 ? T15840 : T15746;
  assign T15746 = T15839 ? T15793 : T15747;
  assign T15747 = T15792 ? T15770 : T15748;
  assign T15748 = T15769 ? T15759 : T15749;
  assign T15749 = T15758 ? twiddle4_2_129_real : twiddle4_2_128_real;
  assign twiddle4_2_128_real = T15752 + T15750;
  assign T15750 = $signed(T15751) / $signed(22'h100000);
  assign T15751 = $signed(31'h2d413ccc) * $signed(16'h0);
  assign T15752 = $signed(T15753) / $signed(22'h100000);
  assign T15753 = $signed(31'h2d413ccc) * $signed(16'h1);
  assign twiddle4_2_129_real = T15756 + T15754;
  assign T15754 = $signed(T15755) / $signed(22'h100000);
  assign T15755 = $signed(31'h2d881ae7) * $signed(16'h0);
  assign T15756 = $signed(T15757) / $signed(22'h100000);
  assign T15757 = $signed(31'h2cf9ef09) * $signed(16'h1);
  assign T15758 = T10817[1'h0:1'h0];
  assign T15759 = T15768 ? twiddle4_2_131_real : twiddle4_2_130_real;
  assign twiddle4_2_130_real = T15762 + T15760;
  assign T15760 = $signed(T15761) / $signed(22'h100000);
  assign T15761 = $signed(31'h2dce88a9) * $signed(16'h0);
  assign T15762 = $signed(T15763) / $signed(22'h100000);
  assign T15763 = $signed(31'h2cb2324b) * $signed(16'h1);
  assign twiddle4_2_131_real = T15766 + T15764;
  assign T15764 = $signed(T15765) / $signed(22'h100000);
  assign T15765 = $signed(31'h2e148566) * $signed(16'h0);
  assign T15766 = $signed(T15767) / $signed(22'h100000);
  assign T15767 = $signed(31'h2c6a0746) * $signed(16'h1);
  assign T15768 = T10817[1'h0:1'h0];
  assign T15769 = T10817[1'h1:1'h1];
  assign T15770 = T15791 ? T15781 : T15771;
  assign T15771 = T15780 ? twiddle4_2_133_real : twiddle4_2_132_real;
  assign twiddle4_2_132_real = T15774 + T15772;
  assign T15772 = $signed(T15773) / $signed(22'h100000);
  assign T15773 = $signed(31'h2e5a106f) * $signed(16'h0);
  assign T15774 = $signed(T15775) / $signed(22'h100000);
  assign T15775 = $signed(31'h2c216eaa) * $signed(16'h1);
  assign twiddle4_2_133_real = T15778 + T15776;
  assign T15776 = $signed(T15777) / $signed(22'h100000);
  assign T15777 = $signed(31'h2e9f291b) * $signed(16'h0);
  assign T15778 = $signed(T15779) / $signed(22'h100000);
  assign T15779 = $signed(31'h2bd8692b) * $signed(16'h1);
  assign T15780 = T10817[1'h0:1'h0];
  assign T15781 = T15790 ? twiddle4_2_135_real : twiddle4_2_134_real;
  assign twiddle4_2_134_real = T15784 + T15782;
  assign T15782 = $signed(T15783) / $signed(22'h100000);
  assign T15783 = $signed(31'h2ee3cebe) * $signed(16'h0);
  assign T15784 = $signed(T15785) / $signed(22'h100000);
  assign T15785 = $signed(31'h2b8ef77c) * $signed(16'h1);
  assign twiddle4_2_135_real = T15788 + T15786;
  assign T15786 = $signed(T15787) / $signed(22'h100000);
  assign T15787 = $signed(31'h2f2800ae) * $signed(16'h0);
  assign T15788 = $signed(T15789) / $signed(22'h100000);
  assign T15789 = $signed(31'h2b451a54) * $signed(16'h1);
  assign T15790 = T10817[1'h0:1'h0];
  assign T15791 = T10817[1'h1:1'h1];
  assign T15792 = T10817[2'h2:2'h2];
  assign T15793 = T15838 ? T15816 : T15794;
  assign T15794 = T15815 ? T15805 : T15795;
  assign T15795 = T15804 ? twiddle4_2_137_real : twiddle4_2_136_real;
  assign twiddle4_2_136_real = T15798 + T15796;
  assign T15796 = $signed(T15797) / $signed(22'h100000);
  assign T15797 = $signed(31'h2f6bbe44) * $signed(16'h0);
  assign T15798 = $signed(T15799) / $signed(22'h100000);
  assign T15799 = $signed(31'h2afad269) * $signed(16'h1);
  assign twiddle4_2_137_real = T15802 + T15800;
  assign T15800 = $signed(T15801) / $signed(22'h100000);
  assign T15801 = $signed(31'h2faf06d9) * $signed(16'h0);
  assign T15802 = $signed(T15803) / $signed(22'h100000);
  assign T15803 = $signed(31'h2ab02071) * $signed(16'h1);
  assign T15804 = T10817[1'h0:1'h0];
  assign T15805 = T15814 ? twiddle4_2_139_real : twiddle4_2_138_real;
  assign twiddle4_2_138_real = T15808 + T15806;
  assign T15806 = $signed(T15807) / $signed(22'h100000);
  assign T15807 = $signed(31'h2ff1d9c6) * $signed(16'h0);
  assign T15808 = $signed(T15809) / $signed(22'h100000);
  assign T15809 = $signed(31'h2a650525) * $signed(16'h1);
  assign twiddle4_2_139_real = T15812 + T15810;
  assign T15810 = $signed(T15811) / $signed(22'h100000);
  assign T15811 = $signed(31'h30343667) * $signed(16'h0);
  assign T15812 = $signed(T15813) / $signed(22'h100000);
  assign T15813 = $signed(31'h2a19813e) * $signed(16'h1);
  assign T15814 = T10817[1'h0:1'h0];
  assign T15815 = T10817[1'h1:1'h1];
  assign T15816 = T15837 ? T15827 : T15817;
  assign T15817 = T15826 ? twiddle4_2_141_real : twiddle4_2_140_real;
  assign twiddle4_2_140_real = T15820 + T15818;
  assign T15818 = $signed(T15819) / $signed(22'h100000);
  assign T15819 = $signed(31'h30761c17) * $signed(16'h0);
  assign T15820 = $signed(T15821) / $signed(22'h100000);
  assign T15821 = $signed(31'h29cd9577) * $signed(16'h1);
  assign twiddle4_2_141_real = T15824 + T15822;
  assign T15822 = $signed(T15823) / $signed(22'h100000);
  assign T15823 = $signed(31'h30b78a35) * $signed(16'h0);
  assign T15824 = $signed(T15825) / $signed(22'h100000);
  assign T15825 = $signed(31'h2981428b) * $signed(16'h1);
  assign T15826 = T10817[1'h0:1'h0];
  assign T15827 = T15836 ? twiddle4_2_143_real : twiddle4_2_142_real;
  assign twiddle4_2_142_real = T15830 + T15828;
  assign T15828 = $signed(T15829) / $signed(22'h100000);
  assign T15829 = $signed(31'h30f8801f) * $signed(16'h0);
  assign T15830 = $signed(T15831) / $signed(22'h100000);
  assign T15831 = $signed(31'h29348937) * $signed(16'h1);
  assign twiddle4_2_143_real = T15834 + T15832;
  assign T15832 = $signed(T15833) / $signed(22'h100000);
  assign T15833 = $signed(31'h3138fd34) * $signed(16'h0);
  assign T15834 = $signed(T15835) / $signed(22'h100000);
  assign T15835 = $signed(31'h28e76a37) * $signed(16'h1);
  assign T15836 = T10817[1'h0:1'h0];
  assign T15837 = T10817[1'h1:1'h1];
  assign T15838 = T10817[2'h2:2'h2];
  assign T15839 = T10817[2'h3:2'h3];
  assign T15840 = T15933 ? T15887 : T15841;
  assign T15841 = T15886 ? T15864 : T15842;
  assign T15842 = T15863 ? T15853 : T15843;
  assign T15843 = T15852 ? twiddle4_2_145_real : twiddle4_2_144_real;
  assign twiddle4_2_144_real = T15846 + T15844;
  assign T15844 = $signed(T15845) / $signed(22'h100000);
  assign T15845 = $signed(31'h317900d6) * $signed(16'h0);
  assign T15846 = $signed(T15847) / $signed(22'h100000);
  assign T15847 = $signed(31'h2899e64a) * $signed(16'h1);
  assign twiddle4_2_145_real = T15850 + T15848;
  assign T15848 = $signed(T15849) / $signed(22'h100000);
  assign T15849 = $signed(31'h31b88a66) * $signed(16'h0);
  assign T15850 = $signed(T15851) / $signed(22'h100000);
  assign T15851 = $signed(31'h284bfe2f) * $signed(16'h1);
  assign T15852 = T10817[1'h0:1'h0];
  assign T15853 = T15862 ? twiddle4_2_147_real : twiddle4_2_146_real;
  assign twiddle4_2_146_real = T15856 + T15854;
  assign T15854 = $signed(T15855) / $signed(22'h100000);
  assign T15855 = $signed(31'h31f79947) * $signed(16'h0);
  assign T15856 = $signed(T15857) / $signed(22'h100000);
  assign T15857 = $signed(31'h27fdb2a6) * $signed(16'h1);
  assign twiddle4_2_147_real = T15860 + T15858;
  assign T15858 = $signed(T15859) / $signed(22'h100000);
  assign T15859 = $signed(31'h32362cdf) * $signed(16'h0);
  assign T15860 = $signed(T15861) / $signed(22'h100000);
  assign T15861 = $signed(31'h27af0471) * $signed(16'h1);
  assign T15862 = T10817[1'h0:1'h0];
  assign T15863 = T10817[1'h1:1'h1];
  assign T15864 = T15885 ? T15875 : T15865;
  assign T15865 = T15874 ? twiddle4_2_149_real : twiddle4_2_148_real;
  assign twiddle4_2_148_real = T15868 + T15866;
  assign T15866 = $signed(T15867) / $signed(22'h100000);
  assign T15867 = $signed(31'h32744493) * $signed(16'h0);
  assign T15868 = $signed(T15869) / $signed(22'h100000);
  assign T15869 = $signed(31'h275ff452) * $signed(16'h1);
  assign twiddle4_2_149_real = T15872 + T15870;
  assign T15870 = $signed(T15871) / $signed(22'h100000);
  assign T15871 = $signed(31'h32b1dfc9) * $signed(16'h0);
  assign T15872 = $signed(T15873) / $signed(22'h100000);
  assign T15873 = $signed(31'h2710830b) * $signed(16'h1);
  assign T15874 = T10817[1'h0:1'h0];
  assign T15875 = T15884 ? twiddle4_2_151_real : twiddle4_2_150_real;
  assign twiddle4_2_150_real = T15878 + T15876;
  assign T15876 = $signed(T15877) / $signed(22'h100000);
  assign T15877 = $signed(31'h32eefde9) * $signed(16'h0);
  assign T15878 = $signed(T15879) / $signed(22'h100000);
  assign T15879 = $signed(31'h26c0b162) * $signed(16'h1);
  assign twiddle4_2_151_real = T15882 + T15880;
  assign T15880 = $signed(T15881) / $signed(22'h100000);
  assign T15881 = $signed(31'h332b9e5d) * $signed(16'h0);
  assign T15882 = $signed(T15883) / $signed(22'h100000);
  assign T15883 = $signed(31'h2670801a) * $signed(16'h1);
  assign T15884 = T10817[1'h0:1'h0];
  assign T15885 = T10817[1'h1:1'h1];
  assign T15886 = T10817[2'h2:2'h2];
  assign T15887 = T15932 ? T15910 : T15888;
  assign T15888 = T15909 ? T15899 : T15889;
  assign T15889 = T15898 ? twiddle4_2_153_real : twiddle4_2_152_real;
  assign twiddle4_2_152_real = T15892 + T15890;
  assign T15890 = $signed(T15891) / $signed(22'h100000);
  assign T15891 = $signed(31'h3367c08f) * $signed(16'h0);
  assign T15892 = $signed(T15893) / $signed(22'h100000);
  assign T15893 = $signed(31'h261feff9) * $signed(16'h1);
  assign twiddle4_2_153_real = T15896 + T15894;
  assign T15894 = $signed(T15895) / $signed(22'h100000);
  assign T15895 = $signed(31'h33a363eb) * $signed(16'h0);
  assign T15896 = $signed(T15897) / $signed(22'h100000);
  assign T15897 = $signed(31'h25cf01c7) * $signed(16'h1);
  assign T15898 = T10817[1'h0:1'h0];
  assign T15899 = T15908 ? twiddle4_2_155_real : twiddle4_2_154_real;
  assign twiddle4_2_154_real = T15902 + T15900;
  assign T15900 = $signed(T15901) / $signed(22'h100000);
  assign T15901 = $signed(31'h33de87de) * $signed(16'h0);
  assign T15902 = $signed(T15903) / $signed(22'h100000);
  assign T15903 = $signed(31'h257db64b) * $signed(16'h1);
  assign twiddle4_2_155_real = T15906 + T15904;
  assign T15904 = $signed(T15905) / $signed(22'h100000);
  assign T15905 = $signed(31'h34192bd5) * $signed(16'h0);
  assign T15906 = $signed(T15907) / $signed(22'h100000);
  assign T15907 = $signed(31'h252c0e4e) * $signed(16'h1);
  assign T15908 = T10817[1'h0:1'h0];
  assign T15909 = T10817[1'h1:1'h1];
  assign T15910 = T15931 ? T15921 : T15911;
  assign T15911 = T15920 ? twiddle4_2_157_real : twiddle4_2_156_real;
  assign twiddle4_2_156_real = T15914 + T15912;
  assign T15912 = $signed(T15913) / $signed(22'h100000);
  assign T15913 = $signed(31'h34534f40) * $signed(16'h0);
  assign T15914 = $signed(T15915) / $signed(22'h100000);
  assign T15915 = $signed(31'h24da0a99) * $signed(16'h1);
  assign twiddle4_2_157_real = T15918 + T15916;
  assign T15916 = $signed(T15917) / $signed(22'h100000);
  assign T15917 = $signed(31'h348cf190) * $signed(16'h0);
  assign T15918 = $signed(T15919) / $signed(22'h100000);
  assign T15919 = $signed(31'h2487abf7) * $signed(16'h1);
  assign T15920 = T10817[1'h0:1'h0];
  assign T15921 = T15930 ? twiddle4_2_159_real : twiddle4_2_158_real;
  assign twiddle4_2_158_real = T15924 + T15922;
  assign T15922 = $signed(T15923) / $signed(22'h100000);
  assign T15923 = $signed(31'h34c61236) * $signed(16'h0);
  assign T15924 = $signed(T15925) / $signed(22'h100000);
  assign T15925 = $signed(31'h2434f332) * $signed(16'h1);
  assign twiddle4_2_159_real = T15928 + T15926;
  assign T15926 = $signed(T15927) / $signed(22'h100000);
  assign T15927 = $signed(31'h34feb0a5) * $signed(16'h0);
  assign T15928 = $signed(T15929) / $signed(22'h100000);
  assign T15929 = $signed(31'h23e1e117) * $signed(16'h1);
  assign T15930 = T10817[1'h0:1'h0];
  assign T15931 = T10817[1'h1:1'h1];
  assign T15932 = T10817[2'h2:2'h2];
  assign T15933 = T10817[2'h3:2'h3];
  assign T15934 = T10817[3'h4:3'h4];
  assign T15935 = T16166 ? T16040 : T15936;
  assign T15936 = T16039 ? T15983 : T15937;
  assign T15937 = T15982 ? T15960 : T15938;
  assign T15938 = T15959 ? T15949 : T15939;
  assign T15939 = T15948 ? twiddle4_2_161_real : twiddle4_2_160_real;
  assign twiddle4_2_160_real = T15942 + T15940;
  assign T15940 = $signed(T15941) / $signed(22'h100000);
  assign T15941 = $signed(31'h3536cc52) * $signed(16'h0);
  assign T15942 = $signed(T15943) / $signed(22'h100000);
  assign T15943 = $signed(31'h238e7673) * $signed(16'h1);
  assign twiddle4_2_161_real = T15946 + T15944;
  assign T15944 = $signed(T15945) / $signed(22'h100000);
  assign T15945 = $signed(31'h356e64b2) * $signed(16'h0);
  assign T15946 = $signed(T15947) / $signed(22'h100000);
  assign T15947 = $signed(31'h233ab413) * $signed(16'h1);
  assign T15948 = T10817[1'h0:1'h0];
  assign T15949 = T15958 ? twiddle4_2_163_real : twiddle4_2_162_real;
  assign twiddle4_2_162_real = T15952 + T15950;
  assign T15950 = $signed(T15951) / $signed(22'h100000);
  assign T15951 = $signed(31'h35a5793c) * $signed(16'h0);
  assign T15952 = $signed(T15953) / $signed(22'h100000);
  assign T15953 = $signed(31'h22e69ac7) * $signed(16'h1);
  assign twiddle4_2_163_real = T15956 + T15954;
  assign T15954 = $signed(T15955) / $signed(22'h100000);
  assign T15955 = $signed(31'h35dc0968) * $signed(16'h0);
  assign T15956 = $signed(T15957) / $signed(22'h100000);
  assign T15957 = $signed(31'h22922b5e) * $signed(16'h1);
  assign T15958 = T10817[1'h0:1'h0];
  assign T15959 = T10817[1'h1:1'h1];
  assign T15960 = T15981 ? T15971 : T15961;
  assign T15961 = T15970 ? twiddle4_2_165_real : twiddle4_2_164_real;
  assign twiddle4_2_164_real = T15964 + T15962;
  assign T15962 = $signed(T15963) / $signed(22'h100000);
  assign T15963 = $signed(31'h361214b0) * $signed(16'h0);
  assign T15964 = $signed(T15965) / $signed(22'h100000);
  assign T15965 = $signed(31'h223d66a8) * $signed(16'h1);
  assign twiddle4_2_165_real = T15968 + T15966;
  assign T15966 = $signed(T15967) / $signed(22'h100000);
  assign T15967 = $signed(31'h36479a8e) * $signed(16'h0);
  assign T15968 = $signed(T15969) / $signed(22'h100000);
  assign T15969 = $signed(31'h21e84d76) * $signed(16'h1);
  assign T15970 = T10817[1'h0:1'h0];
  assign T15971 = T15980 ? twiddle4_2_167_real : twiddle4_2_166_real;
  assign twiddle4_2_166_real = T15974 + T15972;
  assign T15972 = $signed(T15973) / $signed(22'h100000);
  assign T15973 = $signed(31'h367c9a7d) * $signed(16'h0);
  assign T15974 = $signed(T15975) / $signed(22'h100000);
  assign T15975 = $signed(31'h2192e09a) * $signed(16'h1);
  assign twiddle4_2_167_real = T15978 + T15976;
  assign T15976 = $signed(T15977) / $signed(22'h100000);
  assign T15977 = $signed(31'h36b113fd) * $signed(16'h0);
  assign T15978 = $signed(T15979) / $signed(22'h100000);
  assign T15979 = $signed(31'h213d20e8) * $signed(16'h1);
  assign T15980 = T10817[1'h0:1'h0];
  assign T15981 = T10817[1'h1:1'h1];
  assign T15982 = T10817[2'h2:2'h2];
  assign T15983 = T16038 ? T16008 : T15984;
  assign T15984 = T16007 ? T15995 : T15985;
  assign T15985 = T15994 ? twiddle4_2_169_real : twiddle4_2_168_real;
  assign twiddle4_2_168_real = T15988 + T15986;
  assign T15986 = $signed(T15987) / $signed(22'h100000);
  assign T15987 = $signed(31'h36e5068a) * $signed(16'h0);
  assign T15988 = $signed(T15989) / $signed(22'h100000);
  assign T15989 = $signed(31'h20e70f32) * $signed(16'h1);
  assign twiddle4_2_169_real = T15992 + T15990;
  assign T15990 = $signed(T15991) / $signed(22'h100000);
  assign T15991 = $signed(31'h371871a4) * $signed(16'h0);
  assign T15992 = $signed(T15993) / $signed(22'h100000);
  assign T15993 = $signed(31'h2090ac4d) * $signed(16'h1);
  assign T15994 = T10817[1'h0:1'h0];
  assign T15995 = T16006 ? twiddle4_2_171_real : twiddle4_2_170_real;
  assign twiddle4_2_170_real = T15998 + T15996;
  assign T15996 = $signed(T15997) / $signed(22'h100000);
  assign T15997 = $signed(31'h374b54ce) * $signed(16'h0);
  assign T15998 = $signed(T15999) / $signed(22'h100000);
  assign T15999 = $signed(31'h2039f90e) * $signed(16'h1);
  assign twiddle4_2_171_real = T16002 + T16000;
  assign T16000 = $signed(T16001) / $signed(22'h100000);
  assign T16001 = $signed(31'h377daf89) * $signed(16'h0);
  assign T16002 = {T16005, T16003};
  assign T16003 = $signed(T16004) / $signed(22'h100000);
  assign T16004 = $signed(30'h1fe2f64b) * $signed(16'h1);
  assign T16005 = T16003[6'h2d:6'h2d];
  assign T16006 = T10817[1'h0:1'h0];
  assign T16007 = T10817[1'h1:1'h1];
  assign T16008 = T16037 ? T16023 : T16009;
  assign T16009 = T16022 ? twiddle4_2_173_real : twiddle4_2_172_real;
  assign twiddle4_2_172_real = T16012 + T16010;
  assign T16010 = $signed(T16011) / $signed(22'h100000);
  assign T16011 = $signed(31'h37af8158) * $signed(16'h0);
  assign T16012 = {T16015, T16013};
  assign T16013 = $signed(T16014) / $signed(22'h100000);
  assign T16014 = $signed(30'h1f8ba4db) * $signed(16'h1);
  assign T16015 = T16013[6'h2d:6'h2d];
  assign twiddle4_2_173_real = T16018 + T16016;
  assign T16016 = $signed(T16017) / $signed(22'h100000);
  assign T16017 = $signed(31'h37e0c9c2) * $signed(16'h0);
  assign T16018 = {T16021, T16019};
  assign T16019 = $signed(T16020) / $signed(22'h100000);
  assign T16020 = $signed(30'h1f340596) * $signed(16'h1);
  assign T16021 = T16019[6'h2d:6'h2d];
  assign T16022 = T10817[1'h0:1'h0];
  assign T16023 = T16036 ? twiddle4_2_175_real : twiddle4_2_174_real;
  assign twiddle4_2_174_real = T16026 + T16024;
  assign T16024 = $signed(T16025) / $signed(22'h100000);
  assign T16025 = $signed(31'h3811884c) * $signed(16'h0);
  assign T16026 = {T16029, T16027};
  assign T16027 = $signed(T16028) / $signed(22'h100000);
  assign T16028 = $signed(30'h1edc1952) * $signed(16'h1);
  assign T16029 = T16027[6'h2d:6'h2d];
  assign twiddle4_2_175_real = T16032 + T16030;
  assign T16030 = $signed(T16031) / $signed(22'h100000);
  assign T16031 = $signed(31'h3841bc7f) * $signed(16'h0);
  assign T16032 = {T16035, T16033};
  assign T16033 = $signed(T16034) / $signed(22'h100000);
  assign T16034 = $signed(30'h1e83e0ea) * $signed(16'h1);
  assign T16035 = T16033[6'h2d:6'h2d];
  assign T16036 = T10817[1'h0:1'h0];
  assign T16037 = T10817[1'h1:1'h1];
  assign T16038 = T10817[2'h2:2'h2];
  assign T16039 = T10817[2'h3:2'h3];
  assign T16040 = T16165 ? T16103 : T16041;
  assign T16041 = T16102 ? T16072 : T16042;
  assign T16042 = T16071 ? T16057 : T16043;
  assign T16043 = T16056 ? twiddle4_2_177_real : twiddle4_2_176_real;
  assign twiddle4_2_176_real = T16046 + T16044;
  assign T16044 = $signed(T16045) / $signed(22'h100000);
  assign T16045 = $signed(31'h387165e3) * $signed(16'h0);
  assign T16046 = {T16049, T16047};
  assign T16047 = $signed(T16048) / $signed(22'h100000);
  assign T16048 = $signed(30'h1e2b5d38) * $signed(16'h1);
  assign T16049 = T16047[6'h2d:6'h2d];
  assign twiddle4_2_177_real = T16052 + T16050;
  assign T16050 = $signed(T16051) / $signed(22'h100000);
  assign T16051 = $signed(31'h38a08402) * $signed(16'h0);
  assign T16052 = {T16055, T16053};
  assign T16053 = $signed(T16054) / $signed(22'h100000);
  assign T16054 = $signed(30'h1dd28f14) * $signed(16'h1);
  assign T16055 = T16053[6'h2d:6'h2d];
  assign T16056 = T10817[1'h0:1'h0];
  assign T16057 = T16070 ? twiddle4_2_179_real : twiddle4_2_178_real;
  assign twiddle4_2_178_real = T16060 + T16058;
  assign T16058 = $signed(T16059) / $signed(22'h100000);
  assign T16059 = $signed(31'h38cf1669) * $signed(16'h0);
  assign T16060 = {T16063, T16061};
  assign T16061 = $signed(T16062) / $signed(22'h100000);
  assign T16062 = $signed(30'h1d79775b) * $signed(16'h1);
  assign T16063 = T16061[6'h2d:6'h2d];
  assign twiddle4_2_179_real = T16066 + T16064;
  assign T16064 = $signed(T16065) / $signed(22'h100000);
  assign T16065 = $signed(31'h38fd1ca4) * $signed(16'h0);
  assign T16066 = {T16069, T16067};
  assign T16067 = $signed(T16068) / $signed(22'h100000);
  assign T16068 = $signed(30'h1d2016e8) * $signed(16'h1);
  assign T16069 = T16067[6'h2d:6'h2d];
  assign T16070 = T10817[1'h0:1'h0];
  assign T16071 = T10817[1'h1:1'h1];
  assign T16072 = T16101 ? T16087 : T16073;
  assign T16073 = T16086 ? twiddle4_2_181_real : twiddle4_2_180_real;
  assign twiddle4_2_180_real = T16076 + T16074;
  assign T16074 = $signed(T16075) / $signed(22'h100000);
  assign T16075 = $signed(31'h392a9642) * $signed(16'h0);
  assign T16076 = {T16079, T16077};
  assign T16077 = $signed(T16078) / $signed(22'h100000);
  assign T16078 = $signed(30'h1cc66e99) * $signed(16'h1);
  assign T16079 = T16077[6'h2d:6'h2d];
  assign twiddle4_2_181_real = T16082 + T16080;
  assign T16080 = $signed(T16081) / $signed(22'h100000);
  assign T16081 = $signed(31'h395782d3) * $signed(16'h0);
  assign T16082 = {T16085, T16083};
  assign T16083 = $signed(T16084) / $signed(22'h100000);
  assign T16084 = $signed(30'h1c6c7f49) * $signed(16'h1);
  assign T16085 = T16083[6'h2d:6'h2d];
  assign T16086 = T10817[1'h0:1'h0];
  assign T16087 = T16100 ? twiddle4_2_183_real : twiddle4_2_182_real;
  assign twiddle4_2_182_real = T16090 + T16088;
  assign T16088 = $signed(T16089) / $signed(22'h100000);
  assign T16089 = $signed(31'h3983e1e7) * $signed(16'h0);
  assign T16090 = {T16093, T16091};
  assign T16091 = $signed(T16092) / $signed(22'h100000);
  assign T16092 = $signed(30'h1c1249d8) * $signed(16'h1);
  assign T16093 = T16091[6'h2d:6'h2d];
  assign twiddle4_2_183_real = T16096 + T16094;
  assign T16094 = $signed(T16095) / $signed(22'h100000);
  assign T16095 = $signed(31'h39afb313) * $signed(16'h0);
  assign T16096 = {T16099, T16097};
  assign T16097 = $signed(T16098) / $signed(22'h100000);
  assign T16098 = $signed(30'h1bb7cf23) * $signed(16'h1);
  assign T16099 = T16097[6'h2d:6'h2d];
  assign T16100 = T10817[1'h0:1'h0];
  assign T16101 = T10817[1'h1:1'h1];
  assign T16102 = T10817[2'h2:2'h2];
  assign T16103 = T16164 ? T16134 : T16104;
  assign T16104 = T16133 ? T16119 : T16105;
  assign T16105 = T16118 ? twiddle4_2_185_real : twiddle4_2_184_real;
  assign twiddle4_2_184_real = T16108 + T16106;
  assign T16106 = $signed(T16107) / $signed(22'h100000);
  assign T16107 = $signed(31'h39daf5e8) * $signed(16'h0);
  assign T16108 = {T16111, T16109};
  assign T16109 = $signed(T16110) / $signed(22'h100000);
  assign T16110 = $signed(30'h1b5d1009) * $signed(16'h1);
  assign T16111 = T16109[6'h2d:6'h2d];
  assign twiddle4_2_185_real = T16114 + T16112;
  assign T16112 = $signed(T16113) / $signed(22'h100000);
  assign T16113 = $signed(31'h3a05a9fd) * $signed(16'h0);
  assign T16114 = {T16117, T16115};
  assign T16115 = $signed(T16116) / $signed(22'h100000);
  assign T16116 = $signed(30'h1b020d6c) * $signed(16'h1);
  assign T16117 = T16115[6'h2d:6'h2d];
  assign T16118 = T10817[1'h0:1'h0];
  assign T16119 = T16132 ? twiddle4_2_187_real : twiddle4_2_186_real;
  assign twiddle4_2_186_real = T16122 + T16120;
  assign T16120 = $signed(T16121) / $signed(22'h100000);
  assign T16121 = $signed(31'h3a2fcee8) * $signed(16'h0);
  assign T16122 = {T16125, T16123};
  assign T16123 = $signed(T16124) / $signed(22'h100000);
  assign T16124 = $signed(30'h1aa6c82b) * $signed(16'h1);
  assign T16125 = T16123[6'h2d:6'h2d];
  assign twiddle4_2_187_real = T16128 + T16126;
  assign T16126 = $signed(T16127) / $signed(22'h100000);
  assign T16127 = $signed(31'h3a596441) * $signed(16'h0);
  assign T16128 = {T16131, T16129};
  assign T16129 = $signed(T16130) / $signed(22'h100000);
  assign T16130 = $signed(30'h1a4b4127) * $signed(16'h1);
  assign T16131 = T16129[6'h2d:6'h2d];
  assign T16132 = T10817[1'h0:1'h0];
  assign T16133 = T10817[1'h1:1'h1];
  assign T16134 = T16163 ? T16149 : T16135;
  assign T16135 = T16148 ? twiddle4_2_189_real : twiddle4_2_188_real;
  assign twiddle4_2_188_real = T16138 + T16136;
  assign T16136 = $signed(T16137) / $signed(22'h100000);
  assign T16137 = $signed(31'h3a8269a2) * $signed(16'h0);
  assign T16138 = {T16141, T16139};
  assign T16139 = $signed(T16140) / $signed(22'h100000);
  assign T16140 = $signed(30'h19ef7943) * $signed(16'h1);
  assign T16141 = T16139[6'h2d:6'h2d];
  assign twiddle4_2_189_real = T16144 + T16142;
  assign T16142 = $signed(T16143) / $signed(22'h100000);
  assign T16143 = $signed(31'h3aaadea5) * $signed(16'h0);
  assign T16144 = {T16147, T16145};
  assign T16145 = $signed(T16146) / $signed(22'h100000);
  assign T16146 = $signed(30'h19937161) * $signed(16'h1);
  assign T16147 = T16145[6'h2d:6'h2d];
  assign T16148 = T10817[1'h0:1'h0];
  assign T16149 = T16162 ? twiddle4_2_191_real : twiddle4_2_190_real;
  assign twiddle4_2_190_real = T16152 + T16150;
  assign T16150 = $signed(T16151) / $signed(22'h100000);
  assign T16151 = $signed(31'h3ad2c2e7) * $signed(16'h0);
  assign T16152 = {T16155, T16153};
  assign T16153 = $signed(T16154) / $signed(22'h100000);
  assign T16154 = $signed(30'h19372a63) * $signed(16'h1);
  assign T16155 = T16153[6'h2d:6'h2d];
  assign twiddle4_2_191_real = T16158 + T16156;
  assign T16156 = $signed(T16157) / $signed(22'h100000);
  assign T16157 = $signed(31'h3afa1605) * $signed(16'h0);
  assign T16158 = {T16161, T16159};
  assign T16159 = $signed(T16160) / $signed(22'h100000);
  assign T16160 = $signed(30'h18daa52e) * $signed(16'h1);
  assign T16161 = T16159[6'h2d:6'h2d];
  assign T16162 = T10817[1'h0:1'h0];
  assign T16163 = T10817[1'h1:1'h1];
  assign T16164 = T10817[2'h2:2'h2];
  assign T16165 = T10817[2'h3:2'h3];
  assign T16166 = T10817[3'h4:3'h4];
  assign T16167 = T10817[3'h5:3'h5];
  assign T16168 = T16718 ? T16432 : T16169;
  assign T16169 = T16431 ? T16296 : T16170;
  assign T16170 = T16295 ? T16233 : T16171;
  assign T16171 = T16232 ? T16202 : T16172;
  assign T16172 = T16201 ? T16187 : T16173;
  assign T16173 = T16186 ? twiddle4_2_193_real : twiddle4_2_192_real;
  assign twiddle4_2_192_real = T16176 + T16174;
  assign T16174 = $signed(T16175) / $signed(22'h100000);
  assign T16175 = $signed(31'h3b20d79e) * $signed(16'h0);
  assign T16176 = {T16179, T16177};
  assign T16177 = $signed(T16178) / $signed(22'h100000);
  assign T16178 = $signed(30'h187de2a6) * $signed(16'h1);
  assign T16179 = T16177[6'h2d:6'h2d];
  assign twiddle4_2_193_real = T16182 + T16180;
  assign T16180 = $signed(T16181) / $signed(22'h100000);
  assign T16181 = $signed(31'h3b470752) * $signed(16'h0);
  assign T16182 = {T16185, T16183};
  assign T16183 = $signed(T16184) / $signed(22'h100000);
  assign T16184 = $signed(30'h1820e3b0) * $signed(16'h1);
  assign T16185 = T16183[6'h2d:6'h2d];
  assign T16186 = T10817[1'h0:1'h0];
  assign T16187 = T16200 ? twiddle4_2_195_real : twiddle4_2_194_real;
  assign twiddle4_2_194_real = T16190 + T16188;
  assign T16188 = $signed(T16189) / $signed(22'h100000);
  assign T16189 = $signed(31'h3b6ca4c4) * $signed(16'h0);
  assign T16190 = {T16193, T16191};
  assign T16191 = $signed(T16192) / $signed(22'h100000);
  assign T16192 = $signed(30'h17c3a931) * $signed(16'h1);
  assign T16193 = T16191[6'h2d:6'h2d];
  assign twiddle4_2_195_real = T16196 + T16194;
  assign T16194 = $signed(T16195) / $signed(22'h100000);
  assign T16195 = $signed(31'h3b91af96) * $signed(16'h0);
  assign T16196 = {T16199, T16197};
  assign T16197 = $signed(T16198) / $signed(22'h100000);
  assign T16198 = $signed(30'h1766340f) * $signed(16'h1);
  assign T16199 = T16197[6'h2d:6'h2d];
  assign T16200 = T10817[1'h0:1'h0];
  assign T16201 = T10817[1'h1:1'h1];
  assign T16202 = T16231 ? T16217 : T16203;
  assign T16203 = T16216 ? twiddle4_2_197_real : twiddle4_2_196_real;
  assign twiddle4_2_196_real = T16206 + T16204;
  assign T16204 = $signed(T16205) / $signed(22'h100000);
  assign T16205 = $signed(31'h3bb6276d) * $signed(16'h0);
  assign T16206 = {T16209, T16207};
  assign T16207 = $signed(T16208) / $signed(22'h100000);
  assign T16208 = $signed(30'h17088530) * $signed(16'h1);
  assign T16209 = T16207[6'h2d:6'h2d];
  assign twiddle4_2_197_real = T16212 + T16210;
  assign T16210 = $signed(T16211) / $signed(22'h100000);
  assign T16211 = $signed(31'h3bda0bef) * $signed(16'h0);
  assign T16212 = {T16215, T16213};
  assign T16213 = $signed(T16214) / $signed(22'h100000);
  assign T16214 = $signed(30'h16aa9d7d) * $signed(16'h1);
  assign T16215 = T16213[6'h2d:6'h2d];
  assign T16216 = T10817[1'h0:1'h0];
  assign T16217 = T16230 ? twiddle4_2_199_real : twiddle4_2_198_real;
  assign twiddle4_2_198_real = T16220 + T16218;
  assign T16218 = $signed(T16219) / $signed(22'h100000);
  assign T16219 = $signed(31'h3bfd5cc4) * $signed(16'h0);
  assign T16220 = {T16223, T16221};
  assign T16221 = $signed(T16222) / $signed(22'h100000);
  assign T16222 = $signed(30'h164c7ddd) * $signed(16'h1);
  assign T16223 = T16221[6'h2d:6'h2d];
  assign twiddle4_2_199_real = T16226 + T16224;
  assign T16224 = $signed(T16225) / $signed(22'h100000);
  assign T16225 = $signed(31'h3c201994) * $signed(16'h0);
  assign T16226 = {T16229, T16227};
  assign T16227 = $signed(T16228) / $signed(22'h100000);
  assign T16228 = $signed(30'h15ee2737) * $signed(16'h1);
  assign T16229 = T16227[6'h2d:6'h2d];
  assign T16230 = T10817[1'h0:1'h0];
  assign T16231 = T10817[1'h1:1'h1];
  assign T16232 = T10817[2'h2:2'h2];
  assign T16233 = T16294 ? T16264 : T16234;
  assign T16234 = T16263 ? T16249 : T16235;
  assign T16235 = T16248 ? twiddle4_2_201_real : twiddle4_2_200_real;
  assign twiddle4_2_200_real = T16238 + T16236;
  assign T16236 = $signed(T16237) / $signed(22'h100000);
  assign T16237 = $signed(31'h3c424209) * $signed(16'h0);
  assign T16238 = {T16241, T16239};
  assign T16239 = $signed(T16240) / $signed(22'h100000);
  assign T16240 = $signed(30'h158f9a75) * $signed(16'h1);
  assign T16241 = T16239[6'h2d:6'h2d];
  assign twiddle4_2_201_real = T16244 + T16242;
  assign T16242 = $signed(T16243) / $signed(22'h100000);
  assign T16243 = $signed(31'h3c63d5d0) * $signed(16'h0);
  assign T16244 = {T16247, T16245};
  assign T16245 = $signed(T16246) / $signed(22'h100000);
  assign T16246 = $signed(30'h1530d880) * $signed(16'h1);
  assign T16247 = T16245[6'h2d:6'h2d];
  assign T16248 = T10817[1'h0:1'h0];
  assign T16249 = T16262 ? twiddle4_2_203_real : twiddle4_2_202_real;
  assign twiddle4_2_202_real = T16252 + T16250;
  assign T16250 = $signed(T16251) / $signed(22'h100000);
  assign T16251 = $signed(31'h3c84d496) * $signed(16'h0);
  assign T16252 = {T16255, T16253};
  assign T16253 = $signed(T16254) / $signed(22'h100000);
  assign T16254 = $signed(30'h14d1e242) * $signed(16'h1);
  assign T16255 = T16253[6'h2d:6'h2d];
  assign twiddle4_2_203_real = T16258 + T16256;
  assign T16256 = $signed(T16257) / $signed(22'h100000);
  assign T16257 = $signed(31'h3ca53e08) * $signed(16'h0);
  assign T16258 = {T16261, T16259};
  assign T16259 = $signed(T16260) / $signed(22'h100000);
  assign T16260 = $signed(30'h1472b8a5) * $signed(16'h1);
  assign T16261 = T16259[6'h2d:6'h2d];
  assign T16262 = T10817[1'h0:1'h0];
  assign T16263 = T10817[1'h1:1'h1];
  assign T16264 = T16293 ? T16279 : T16265;
  assign T16265 = T16278 ? twiddle4_2_205_real : twiddle4_2_204_real;
  assign twiddle4_2_204_real = T16268 + T16266;
  assign T16266 = $signed(T16267) / $signed(22'h100000);
  assign T16267 = $signed(31'h3cc511d8) * $signed(16'h0);
  assign T16268 = {T16271, T16269};
  assign T16269 = $signed(T16270) / $signed(22'h100000);
  assign T16270 = $signed(30'h14135c94) * $signed(16'h1);
  assign T16271 = T16269[6'h2d:6'h2d];
  assign twiddle4_2_205_real = T16274 + T16272;
  assign T16272 = $signed(T16273) / $signed(22'h100000);
  assign T16273 = $signed(31'h3ce44fb6) * $signed(16'h0);
  assign T16274 = {T16277, T16275};
  assign T16275 = $signed(T16276) / $signed(22'h100000);
  assign T16276 = $signed(30'h13b3cefa) * $signed(16'h1);
  assign T16277 = T16275[6'h2d:6'h2d];
  assign T16278 = T10817[1'h0:1'h0];
  assign T16279 = T16292 ? twiddle4_2_207_real : twiddle4_2_206_real;
  assign twiddle4_2_206_real = T16282 + T16280;
  assign T16280 = $signed(T16281) / $signed(22'h100000);
  assign T16281 = $signed(31'h3d02f756) * $signed(16'h0);
  assign T16282 = {T16285, T16283};
  assign T16283 = $signed(T16284) / $signed(22'h100000);
  assign T16284 = $signed(30'h135410c2) * $signed(16'h1);
  assign T16285 = T16283[6'h2d:6'h2d];
  assign twiddle4_2_207_real = T16288 + T16286;
  assign T16286 = $signed(T16287) / $signed(22'h100000);
  assign T16287 = $signed(31'h3d21086c) * $signed(16'h0);
  assign T16288 = {T16291, T16289};
  assign T16289 = $signed(T16290) / $signed(22'h100000);
  assign T16290 = $signed(30'h12f422da) * $signed(16'h1);
  assign T16291 = T16289[6'h2d:6'h2d];
  assign T16292 = T10817[1'h0:1'h0];
  assign T16293 = T10817[1'h1:1'h1];
  assign T16294 = T10817[2'h2:2'h2];
  assign T16295 = T10817[2'h3:2'h3];
  assign T16296 = T16430 ? T16360 : T16297;
  assign T16297 = T16359 ? T16328 : T16298;
  assign T16298 = T16327 ? T16313 : T16299;
  assign T16299 = T16312 ? twiddle4_2_209_real : twiddle4_2_208_real;
  assign twiddle4_2_208_real = T16302 + T16300;
  assign T16300 = $signed(T16301) / $signed(22'h100000);
  assign T16301 = $signed(31'h3d3e82ad) * $signed(16'h0);
  assign T16302 = {T16305, T16303};
  assign T16303 = $signed(T16304) / $signed(22'h100000);
  assign T16304 = $signed(30'h1294062e) * $signed(16'h1);
  assign T16305 = T16303[6'h2d:6'h2d];
  assign twiddle4_2_209_real = T16308 + T16306;
  assign T16306 = $signed(T16307) / $signed(22'h100000);
  assign T16307 = $signed(31'h3d5b65d1) * $signed(16'h0);
  assign T16308 = {T16311, T16309};
  assign T16309 = $signed(T16310) / $signed(22'h100000);
  assign T16310 = $signed(30'h1233bbab) * $signed(16'h1);
  assign T16311 = T16309[6'h2d:6'h2d];
  assign T16312 = T10817[1'h0:1'h0];
  assign T16313 = T16326 ? twiddle4_2_211_real : twiddle4_2_210_real;
  assign twiddle4_2_210_real = T16316 + T16314;
  assign T16314 = $signed(T16315) / $signed(22'h100000);
  assign T16315 = $signed(31'h3d77b191) * $signed(16'h0);
  assign T16316 = {T16319, T16317};
  assign T16317 = $signed(T16318) / $signed(22'h100000);
  assign T16318 = $signed(30'h11d3443f) * $signed(16'h1);
  assign T16319 = T16317[6'h2d:6'h2d];
  assign twiddle4_2_211_real = T16322 + T16320;
  assign T16320 = $signed(T16321) / $signed(22'h100000);
  assign T16321 = $signed(31'h3d9365a7) * $signed(16'h0);
  assign T16322 = {T16325, T16323};
  assign T16323 = $signed(T16324) / $signed(22'h100000);
  assign T16324 = $signed(30'h1172a0d7) * $signed(16'h1);
  assign T16325 = T16323[6'h2d:6'h2d];
  assign T16326 = T10817[1'h0:1'h0];
  assign T16327 = T10817[1'h1:1'h1];
  assign T16328 = T16358 ? T16343 : T16329;
  assign T16329 = T16342 ? twiddle4_2_213_real : twiddle4_2_212_real;
  assign twiddle4_2_212_real = T16332 + T16330;
  assign T16330 = $signed(T16331) / $signed(22'h100000);
  assign T16331 = $signed(31'h3dae81ce) * $signed(16'h0);
  assign T16332 = {T16335, T16333};
  assign T16333 = $signed(T16334) / $signed(22'h100000);
  assign T16334 = $signed(30'h1111d262) * $signed(16'h1);
  assign T16335 = T16333[6'h2d:6'h2d];
  assign twiddle4_2_213_real = T16338 + T16336;
  assign T16336 = $signed(T16337) / $signed(22'h100000);
  assign T16337 = $signed(31'h3dc905c4) * $signed(16'h0);
  assign T16338 = {T16341, T16339};
  assign T16339 = $signed(T16340) / $signed(22'h100000);
  assign T16340 = $signed(30'h10b0d9cf) * $signed(16'h1);
  assign T16341 = T16339[6'h2d:6'h2d];
  assign T16342 = T10817[1'h0:1'h0];
  assign T16343 = T16357 ? twiddle4_2_215_real : twiddle4_2_214_real;
  assign twiddle4_2_214_real = T16346 + T16344;
  assign T16344 = $signed(T16345) / $signed(22'h100000);
  assign T16345 = $signed(31'h3de2f147) * $signed(16'h0);
  assign T16346 = {T16349, T16347};
  assign T16347 = $signed(T16348) / $signed(22'h100000);
  assign T16348 = $signed(30'h104fb80e) * $signed(16'h1);
  assign T16349 = T16347[6'h2d:6'h2d];
  assign twiddle4_2_215_real = T16352 + T16350;
  assign T16350 = $signed(T16351) / $signed(22'h100000);
  assign T16351 = $signed(31'h3dfc4418) * $signed(16'h0);
  assign T16352 = {T16355, T16353};
  assign T16353 = $signed(T16354) / $signed(22'h100000);
  assign T16354 = $signed(29'hfee6e0d) * $signed(16'h1);
  assign T16355 = T16356 ? 2'h3 : 2'h0;
  assign T16356 = T16353[6'h2c:6'h2c];
  assign T16357 = T10817[1'h0:1'h0];
  assign T16358 = T10817[1'h1:1'h1];
  assign T16359 = T10817[2'h2:2'h2];
  assign T16360 = T16429 ? T16395 : T16361;
  assign T16361 = T16394 ? T16378 : T16362;
  assign T16362 = T16377 ? twiddle4_2_217_real : twiddle4_2_216_real;
  assign twiddle4_2_216_real = T16365 + T16363;
  assign T16363 = $signed(T16364) / $signed(22'h100000);
  assign T16364 = $signed(31'h3e14fdf7) * $signed(16'h0);
  assign T16365 = {T16368, T16366};
  assign T16366 = $signed(T16367) / $signed(22'h100000);
  assign T16367 = $signed(29'hf8cfcbd) * $signed(16'h1);
  assign T16368 = T16369 ? 2'h3 : 2'h0;
  assign T16369 = T16366[6'h2c:6'h2c];
  assign twiddle4_2_217_real = T16372 + T16370;
  assign T16370 = $signed(T16371) / $signed(22'h100000);
  assign T16371 = $signed(31'h3e2d1ea7) * $signed(16'h0);
  assign T16372 = {T16375, T16373};
  assign T16373 = $signed(T16374) / $signed(22'h100000);
  assign T16374 = $signed(29'hf2b650f) * $signed(16'h1);
  assign T16375 = T16376 ? 2'h3 : 2'h0;
  assign T16376 = T16373[6'h2c:6'h2c];
  assign T16377 = T10817[1'h0:1'h0];
  assign T16378 = T16393 ? twiddle4_2_219_real : twiddle4_2_218_real;
  assign twiddle4_2_218_real = T16381 + T16379;
  assign T16379 = $signed(T16380) / $signed(22'h100000);
  assign T16380 = $signed(31'h3e44a5ee) * $signed(16'h0);
  assign T16381 = {T16384, T16382};
  assign T16382 = $signed(T16383) / $signed(22'h100000);
  assign T16383 = $signed(29'hec9a7f2) * $signed(16'h1);
  assign T16384 = T16385 ? 2'h3 : 2'h0;
  assign T16385 = T16382[6'h2c:6'h2c];
  assign twiddle4_2_219_real = T16388 + T16386;
  assign T16386 = $signed(T16387) / $signed(22'h100000);
  assign T16387 = $signed(31'h3e5b9392) * $signed(16'h0);
  assign T16388 = {T16391, T16389};
  assign T16389 = $signed(T16390) / $signed(22'h100000);
  assign T16390 = $signed(29'he67c659) * $signed(16'h1);
  assign T16391 = T16392 ? 2'h3 : 2'h0;
  assign T16392 = T16389[6'h2c:6'h2c];
  assign T16393 = T10817[1'h0:1'h0];
  assign T16394 = T10817[1'h1:1'h1];
  assign T16395 = T16428 ? T16412 : T16396;
  assign T16396 = T16411 ? twiddle4_2_221_real : twiddle4_2_220_real;
  assign twiddle4_2_220_real = T16399 + T16397;
  assign T16397 = $signed(T16398) / $signed(22'h100000);
  assign T16398 = $signed(31'h3e71e758) * $signed(16'h0);
  assign T16399 = {T16402, T16400};
  assign T16400 = $signed(T16401) / $signed(22'h100000);
  assign T16401 = $signed(29'he05c135) * $signed(16'h1);
  assign T16402 = T16403 ? 2'h3 : 2'h0;
  assign T16403 = T16400[6'h2c:6'h2c];
  assign twiddle4_2_221_real = T16406 + T16404;
  assign T16404 = $signed(T16405) / $signed(22'h100000);
  assign T16405 = $signed(31'h3e87a10b) * $signed(16'h0);
  assign T16406 = {T16409, T16407};
  assign T16407 = $signed(T16408) / $signed(22'h100000);
  assign T16408 = $signed(29'hda39977) * $signed(16'h1);
  assign T16409 = T16410 ? 2'h3 : 2'h0;
  assign T16410 = T16407[6'h2c:6'h2c];
  assign T16411 = T10817[1'h0:1'h0];
  assign T16412 = T16427 ? twiddle4_2_223_real : twiddle4_2_222_real;
  assign twiddle4_2_222_real = T16415 + T16413;
  assign T16413 = $signed(T16414) / $signed(22'h100000);
  assign T16414 = $signed(31'h3e9cc076) * $signed(16'h0);
  assign T16415 = {T16418, T16416};
  assign T16416 = $signed(T16417) / $signed(22'h100000);
  assign T16417 = $signed(29'hd415012) * $signed(16'h1);
  assign T16418 = T16419 ? 2'h3 : 2'h0;
  assign T16419 = T16416[6'h2c:6'h2c];
  assign twiddle4_2_223_real = T16422 + T16420;
  assign T16420 = $signed(T16421) / $signed(22'h100000);
  assign T16421 = $signed(31'h3eb14562) * $signed(16'h0);
  assign T16422 = {T16425, T16423};
  assign T16423 = $signed(T16424) / $signed(22'h100000);
  assign T16424 = $signed(29'hcdee5f9) * $signed(16'h1);
  assign T16425 = T16426 ? 2'h3 : 2'h0;
  assign T16426 = T16423[6'h2c:6'h2c];
  assign T16427 = T10817[1'h0:1'h0];
  assign T16428 = T10817[1'h1:1'h1];
  assign T16429 = T10817[2'h2:2'h2];
  assign T16430 = T10817[2'h3:2'h3];
  assign T16431 = T10817[3'h4:3'h4];
  assign T16432 = T16717 ? T16575 : T16433;
  assign T16433 = T16574 ? T16504 : T16434;
  assign T16434 = T16503 ? T16469 : T16435;
  assign T16435 = T16468 ? T16452 : T16436;
  assign T16436 = T16451 ? twiddle4_2_225_real : twiddle4_2_224_real;
  assign twiddle4_2_224_real = T16439 + T16437;
  assign T16437 = $signed(T16438) / $signed(22'h100000);
  assign T16438 = $signed(31'h3ec52f9f) * $signed(16'h0);
  assign T16439 = {T16442, T16440};
  assign T16440 = $signed(T16441) / $signed(22'h100000);
  assign T16441 = $signed(29'hc7c5c1e) * $signed(16'h1);
  assign T16442 = T16443 ? 2'h3 : 2'h0;
  assign T16443 = T16440[6'h2c:6'h2c];
  assign twiddle4_2_225_real = T16446 + T16444;
  assign T16444 = $signed(T16445) / $signed(22'h100000);
  assign T16445 = $signed(31'h3ed87efb) * $signed(16'h0);
  assign T16446 = {T16449, T16447};
  assign T16447 = $signed(T16448) / $signed(22'h100000);
  assign T16448 = $signed(29'hc19b374) * $signed(16'h1);
  assign T16449 = T16450 ? 2'h3 : 2'h0;
  assign T16450 = T16447[6'h2c:6'h2c];
  assign T16451 = T10817[1'h0:1'h0];
  assign T16452 = T16467 ? twiddle4_2_227_real : twiddle4_2_226_real;
  assign twiddle4_2_226_real = T16455 + T16453;
  assign T16453 = $signed(T16454) / $signed(22'h100000);
  assign T16454 = $signed(31'h3eeb3347) * $signed(16'h0);
  assign T16455 = {T16458, T16456};
  assign T16456 = $signed(T16457) / $signed(22'h100000);
  assign T16457 = $signed(29'hbb6ecef) * $signed(16'h1);
  assign T16458 = T16459 ? 2'h3 : 2'h0;
  assign T16459 = T16456[6'h2c:6'h2c];
  assign twiddle4_2_227_real = T16462 + T16460;
  assign T16460 = $signed(T16461) / $signed(22'h100000);
  assign T16461 = $signed(31'h3efd4c53) * $signed(16'h0);
  assign T16462 = {T16465, T16463};
  assign T16463 = $signed(T16464) / $signed(22'h100000);
  assign T16464 = $signed(29'hb540982) * $signed(16'h1);
  assign T16465 = T16466 ? 2'h3 : 2'h0;
  assign T16466 = T16463[6'h2c:6'h2c];
  assign T16467 = T10817[1'h0:1'h0];
  assign T16468 = T10817[1'h1:1'h1];
  assign T16469 = T16502 ? T16486 : T16470;
  assign T16470 = T16485 ? twiddle4_2_229_real : twiddle4_2_228_real;
  assign twiddle4_2_228_real = T16473 + T16471;
  assign T16471 = $signed(T16472) / $signed(22'h100000);
  assign T16472 = $signed(31'h3f0ec9f4) * $signed(16'h0);
  assign T16473 = {T16476, T16474};
  assign T16474 = $signed(T16475) / $signed(22'h100000);
  assign T16475 = $signed(29'haf10a22) * $signed(16'h1);
  assign T16476 = T16477 ? 2'h3 : 2'h0;
  assign T16477 = T16474[6'h2c:6'h2c];
  assign twiddle4_2_229_real = T16480 + T16478;
  assign T16478 = $signed(T16479) / $signed(22'h100000);
  assign T16479 = $signed(31'h3f1fabff) * $signed(16'h0);
  assign T16480 = {T16483, T16481};
  assign T16481 = $signed(T16482) / $signed(22'h100000);
  assign T16482 = $signed(29'ha8defc2) * $signed(16'h1);
  assign T16483 = T16484 ? 2'h3 : 2'h0;
  assign T16484 = T16481[6'h2c:6'h2c];
  assign T16485 = T10817[1'h0:1'h0];
  assign T16486 = T16501 ? twiddle4_2_231_real : twiddle4_2_230_real;
  assign twiddle4_2_230_real = T16489 + T16487;
  assign T16487 = $signed(T16488) / $signed(22'h100000);
  assign T16488 = $signed(31'h3f2ff249) * $signed(16'h0);
  assign T16489 = {T16492, T16490};
  assign T16490 = $signed(T16491) / $signed(22'h100000);
  assign T16491 = $signed(29'ha2abb58) * $signed(16'h1);
  assign T16492 = T16493 ? 2'h3 : 2'h0;
  assign T16493 = T16490[6'h2c:6'h2c];
  assign twiddle4_2_231_real = T16496 + T16494;
  assign T16494 = $signed(T16495) / $signed(22'h100000);
  assign T16495 = $signed(31'h3f3f9cab) * $signed(16'h0);
  assign T16496 = {T16499, T16497};
  assign T16497 = $signed(T16498) / $signed(22'h100000);
  assign T16498 = $signed(29'h9c76dd8) * $signed(16'h1);
  assign T16499 = T16500 ? 2'h3 : 2'h0;
  assign T16500 = T16497[6'h2c:6'h2c];
  assign T16501 = T10817[1'h0:1'h0];
  assign T16502 = T10817[1'h1:1'h1];
  assign T16503 = T10817[2'h2:2'h2];
  assign T16504 = T16573 ? T16539 : T16505;
  assign T16505 = T16538 ? T16522 : T16506;
  assign T16506 = T16521 ? twiddle4_2_233_real : twiddle4_2_232_real;
  assign twiddle4_2_232_real = T16509 + T16507;
  assign T16507 = $signed(T16508) / $signed(22'h100000);
  assign T16508 = $signed(31'h3f4eaafe) * $signed(16'h0);
  assign T16509 = {T16512, T16510};
  assign T16510 = $signed(T16511) / $signed(22'h100000);
  assign T16511 = $signed(29'h9640837) * $signed(16'h1);
  assign T16512 = T16513 ? 2'h3 : 2'h0;
  assign T16513 = T16510[6'h2c:6'h2c];
  assign twiddle4_2_233_real = T16516 + T16514;
  assign T16514 = $signed(T16515) / $signed(22'h100000);
  assign T16515 = $signed(31'h3f5d1d1c) * $signed(16'h0);
  assign T16516 = {T16519, T16517};
  assign T16517 = $signed(T16518) / $signed(22'h100000);
  assign T16518 = $signed(29'h9008b6a) * $signed(16'h1);
  assign T16519 = T16520 ? 2'h3 : 2'h0;
  assign T16520 = T16517[6'h2c:6'h2c];
  assign T16521 = T10817[1'h0:1'h0];
  assign T16522 = T16537 ? twiddle4_2_235_real : twiddle4_2_234_real;
  assign twiddle4_2_234_real = T16525 + T16523;
  assign T16523 = $signed(T16524) / $signed(22'h100000);
  assign T16524 = $signed(31'h3f6af2e3) * $signed(16'h0);
  assign T16525 = {T16528, T16526};
  assign T16526 = $signed(T16527) / $signed(22'h100000);
  assign T16527 = $signed(29'h89cf867) * $signed(16'h1);
  assign T16528 = T16529 ? 2'h3 : 2'h0;
  assign T16529 = T16526[6'h2c:6'h2c];
  assign twiddle4_2_235_real = T16532 + T16530;
  assign T16530 = $signed(T16531) / $signed(22'h100000);
  assign T16531 = $signed(31'h3f782c2f) * $signed(16'h0);
  assign T16532 = {T16535, T16533};
  assign T16533 = $signed(T16534) / $signed(22'h100000);
  assign T16534 = $signed(29'h8395023) * $signed(16'h1);
  assign T16535 = T16536 ? 2'h3 : 2'h0;
  assign T16536 = T16533[6'h2c:6'h2c];
  assign T16537 = T10817[1'h0:1'h0];
  assign T16538 = T10817[1'h1:1'h1];
  assign T16539 = T16572 ? T16556 : T16540;
  assign T16540 = T16555 ? twiddle4_2_237_real : twiddle4_2_236_real;
  assign twiddle4_2_236_real = T16543 + T16541;
  assign T16541 = $signed(T16542) / $signed(22'h100000);
  assign T16542 = $signed(31'h3f84c8e1) * $signed(16'h0);
  assign T16543 = {T16546, T16544};
  assign T16544 = $signed(T16545) / $signed(22'h100000);
  assign T16545 = $signed(28'h7d59395) * $signed(16'h1);
  assign T16546 = T16547 ? 3'h7 : 3'h0;
  assign T16547 = T16544[6'h2b:6'h2b];
  assign twiddle4_2_237_real = T16550 + T16548;
  assign T16548 = $signed(T16549) / $signed(22'h100000);
  assign T16549 = $signed(31'h3f90c8d9) * $signed(16'h0);
  assign T16550 = {T16553, T16551};
  assign T16551 = $signed(T16552) / $signed(22'h100000);
  assign T16552 = $signed(28'h771c3b2) * $signed(16'h1);
  assign T16553 = T16554 ? 3'h7 : 3'h0;
  assign T16554 = T16551[6'h2b:6'h2b];
  assign T16555 = T10817[1'h0:1'h0];
  assign T16556 = T16571 ? twiddle4_2_239_real : twiddle4_2_238_real;
  assign twiddle4_2_238_real = T16559 + T16557;
  assign T16557 = $signed(T16558) / $signed(22'h100000);
  assign T16558 = $signed(31'h3f9c2bfa) * $signed(16'h0);
  assign T16559 = {T16562, T16560};
  assign T16560 = $signed(T16561) / $signed(22'h100000);
  assign T16561 = $signed(28'h70de171) * $signed(16'h1);
  assign T16562 = T16563 ? 3'h7 : 3'h0;
  assign T16563 = T16560[6'h2b:6'h2b];
  assign twiddle4_2_239_real = T16566 + T16564;
  assign T16564 = $signed(T16565) / $signed(22'h100000);
  assign T16565 = $signed(31'h3fa6f228) * $signed(16'h0);
  assign T16566 = {T16569, T16567};
  assign T16567 = $signed(T16568) / $signed(22'h100000);
  assign T16568 = $signed(28'h6a9edc9) * $signed(16'h1);
  assign T16569 = T16570 ? 3'h7 : 3'h0;
  assign T16570 = T16567[6'h2b:6'h2b];
  assign T16571 = T10817[1'h0:1'h0];
  assign T16572 = T10817[1'h1:1'h1];
  assign T16573 = T10817[2'h2:2'h2];
  assign T16574 = T10817[2'h3:2'h3];
  assign T16575 = T16716 ? T16646 : T16576;
  assign T16576 = T16645 ? T16611 : T16577;
  assign T16577 = T16610 ? T16594 : T16578;
  assign T16578 = T16593 ? twiddle4_2_241_real : twiddle4_2_240_real;
  assign twiddle4_2_240_real = T16581 + T16579;
  assign T16579 = $signed(T16580) / $signed(22'h100000);
  assign T16580 = $signed(31'h3fb11b47) * $signed(16'h0);
  assign T16581 = {T16584, T16582};
  assign T16582 = $signed(T16583) / $signed(22'h100000);
  assign T16583 = $signed(28'h645e9af) * $signed(16'h1);
  assign T16584 = T16585 ? 3'h7 : 3'h0;
  assign T16585 = T16582[6'h2b:6'h2b];
  assign twiddle4_2_241_real = T16588 + T16586;
  assign T16586 = $signed(T16587) / $signed(22'h100000);
  assign T16587 = $signed(31'h3fbaa73f) * $signed(16'h0);
  assign T16588 = {T16591, T16589};
  assign T16589 = $signed(T16590) / $signed(22'h100000);
  assign T16590 = $signed(28'h5e1d61a) * $signed(16'h1);
  assign T16591 = T16592 ? 3'h7 : 3'h0;
  assign T16592 = T16589[6'h2b:6'h2b];
  assign T16593 = T10817[1'h0:1'h0];
  assign T16594 = T16609 ? twiddle4_2_243_real : twiddle4_2_242_real;
  assign twiddle4_2_242_real = T16597 + T16595;
  assign T16595 = $signed(T16596) / $signed(22'h100000);
  assign T16596 = $signed(31'h3fc395f9) * $signed(16'h0);
  assign T16597 = {T16600, T16598};
  assign T16598 = $signed(T16599) / $signed(22'h100000);
  assign T16599 = $signed(28'h57db402) * $signed(16'h1);
  assign T16600 = T16601 ? 3'h7 : 3'h0;
  assign T16601 = T16598[6'h2b:6'h2b];
  assign twiddle4_2_243_real = T16604 + T16602;
  assign T16602 = $signed(T16603) / $signed(22'h100000);
  assign T16603 = $signed(31'h3fcbe75e) * $signed(16'h0);
  assign T16604 = {T16607, T16605};
  assign T16605 = $signed(T16606) / $signed(22'h100000);
  assign T16606 = $signed(28'h519845e) * $signed(16'h1);
  assign T16607 = T16608 ? 3'h7 : 3'h0;
  assign T16608 = T16605[6'h2b:6'h2b];
  assign T16609 = T10817[1'h0:1'h0];
  assign T16610 = T10817[1'h1:1'h1];
  assign T16611 = T16644 ? T16628 : T16612;
  assign T16612 = T16627 ? twiddle4_2_245_real : twiddle4_2_244_real;
  assign twiddle4_2_244_real = T16615 + T16613;
  assign T16613 = $signed(T16614) / $signed(22'h100000);
  assign T16614 = $signed(31'h3fd39b5a) * $signed(16'h0);
  assign T16615 = {T16618, T16616};
  assign T16616 = $signed(T16617) / $signed(22'h100000);
  assign T16617 = $signed(28'h4b54824) * $signed(16'h1);
  assign T16618 = T16619 ? 3'h7 : 3'h0;
  assign T16619 = T16616[6'h2b:6'h2b];
  assign twiddle4_2_245_real = T16622 + T16620;
  assign T16620 = $signed(T16621) / $signed(22'h100000);
  assign T16621 = $signed(31'h3fdab1d9) * $signed(16'h0);
  assign T16622 = {T16625, T16623};
  assign T16623 = $signed(T16624) / $signed(22'h100000);
  assign T16624 = $signed(28'h451004d) * $signed(16'h1);
  assign T16625 = T16626 ? 3'h7 : 3'h0;
  assign T16626 = T16623[6'h2b:6'h2b];
  assign T16627 = T10817[1'h0:1'h0];
  assign T16628 = T16643 ? twiddle4_2_247_real : twiddle4_2_246_real;
  assign twiddle4_2_246_real = T16631 + T16629;
  assign T16629 = $signed(T16630) / $signed(22'h100000);
  assign T16630 = $signed(31'h3fe12acb) * $signed(16'h0);
  assign T16631 = {T16634, T16632};
  assign T16632 = $signed(T16633) / $signed(22'h100000);
  assign T16633 = $signed(27'h3ecadcf) * $signed(16'h1);
  assign T16634 = T16635 ? 4'hf : 4'h0;
  assign T16635 = T16632[6'h2a:6'h2a];
  assign twiddle4_2_247_real = T16638 + T16636;
  assign T16636 = $signed(T16637) / $signed(22'h100000);
  assign T16637 = $signed(31'h3fe7061f) * $signed(16'h0);
  assign T16638 = {T16641, T16639};
  assign T16639 = $signed(T16640) / $signed(22'h100000);
  assign T16640 = $signed(27'h38851a2) * $signed(16'h1);
  assign T16641 = T16642 ? 4'hf : 4'h0;
  assign T16642 = T16639[6'h2a:6'h2a];
  assign T16643 = T10817[1'h0:1'h0];
  assign T16644 = T10817[1'h1:1'h1];
  assign T16645 = T10817[2'h2:2'h2];
  assign T16646 = T16715 ? T16681 : T16647;
  assign T16647 = T16680 ? T16664 : T16648;
  assign T16648 = T16663 ? twiddle4_2_249_real : twiddle4_2_248_real;
  assign twiddle4_2_248_real = T16651 + T16649;
  assign T16649 = $signed(T16650) / $signed(22'h100000);
  assign T16650 = $signed(31'h3fec43c6) * $signed(16'h0);
  assign T16651 = {T16654, T16652};
  assign T16652 = $signed(T16653) / $signed(22'h100000);
  assign T16653 = $signed(27'h323ecbe) * $signed(16'h1);
  assign T16654 = T16655 ? 4'hf : 4'h0;
  assign T16655 = T16652[6'h2a:6'h2a];
  assign twiddle4_2_249_real = T16658 + T16656;
  assign T16656 = $signed(T16657) / $signed(22'h100000);
  assign T16657 = $signed(31'h3ff0e3b5) * $signed(16'h0);
  assign T16658 = {T16661, T16659};
  assign T16659 = $signed(T16660) / $signed(22'h100000);
  assign T16660 = $signed(27'h2bf801a) * $signed(16'h1);
  assign T16661 = T16662 ? 4'hf : 4'h0;
  assign T16662 = T16659[6'h2a:6'h2a];
  assign T16663 = T10817[1'h0:1'h0];
  assign T16664 = T16679 ? twiddle4_2_251_real : twiddle4_2_250_real;
  assign twiddle4_2_250_real = T16667 + T16665;
  assign T16665 = $signed(T16666) / $signed(22'h100000);
  assign T16666 = $signed(31'h3ff4e5df) * $signed(16'h0);
  assign T16667 = {T16670, T16668};
  assign T16668 = $signed(T16669) / $signed(22'h100000);
  assign T16669 = $signed(27'h25b0cae) * $signed(16'h1);
  assign T16670 = T16671 ? 4'hf : 4'h0;
  assign T16671 = T16668[6'h2a:6'h2a];
  assign twiddle4_2_251_real = T16674 + T16672;
  assign T16672 = $signed(T16673) / $signed(22'h100000);
  assign T16673 = $signed(31'h3ff84a3b) * $signed(16'h0);
  assign T16674 = {T16677, T16675};
  assign T16675 = $signed(T16676) / $signed(22'h100000);
  assign T16676 = $signed(26'h1f69373) * $signed(16'h1);
  assign T16677 = T16678 ? 5'h1f : 5'h0;
  assign T16678 = T16675[6'h29:6'h29];
  assign T16679 = T10817[1'h0:1'h0];
  assign T16680 = T10817[1'h1:1'h1];
  assign T16681 = T16714 ? T16698 : T16682;
  assign T16682 = T16697 ? twiddle4_2_253_real : twiddle4_2_252_real;
  assign twiddle4_2_252_real = T16685 + T16683;
  assign T16683 = $signed(T16684) / $signed(22'h100000);
  assign T16684 = $signed(31'h3ffb10c1) * $signed(16'h0);
  assign T16685 = {T16688, T16686};
  assign T16686 = $signed(T16687) / $signed(22'h100000);
  assign T16687 = $signed(26'h192155f) * $signed(16'h1);
  assign T16688 = T16689 ? 5'h1f : 5'h0;
  assign T16689 = T16686[6'h29:6'h29];
  assign twiddle4_2_253_real = T16692 + T16690;
  assign T16690 = $signed(T16691) / $signed(22'h100000);
  assign T16691 = $signed(31'h3ffd3968) * $signed(16'h0);
  assign T16692 = {T16695, T16693};
  assign T16693 = $signed(T16694) / $signed(22'h100000);
  assign T16694 = $signed(26'h12d936b) * $signed(16'h1);
  assign T16695 = T16696 ? 5'h1f : 5'h0;
  assign T16696 = T16693[6'h29:6'h29];
  assign T16697 = T10817[1'h0:1'h0];
  assign T16698 = T16713 ? twiddle4_2_255_real : twiddle4_2_254_real;
  assign twiddle4_2_254_real = T16701 + T16699;
  assign T16699 = $signed(T16700) / $signed(22'h100000);
  assign T16700 = $signed(31'h3ffec42d) * $signed(16'h0);
  assign T16701 = {T16704, T16702};
  assign T16702 = $signed(T16703) / $signed(22'h100000);
  assign T16703 = $signed(25'hc90e8f) * $signed(16'h1);
  assign T16704 = T16705 ? 6'h3f : 6'h0;
  assign T16705 = T16702[6'h28:6'h28];
  assign twiddle4_2_255_real = T16708 + T16706;
  assign T16706 = $signed(T16707) / $signed(22'h100000);
  assign T16707 = $signed(31'h3fffb10b) * $signed(16'h0);
  assign T16708 = {T16711, T16709};
  assign T16709 = $signed(T16710) / $signed(22'h100000);
  assign T16710 = $signed(24'h6487c3) * $signed(16'h1);
  assign T16711 = T16712 ? 7'h7f : 7'h0;
  assign T16712 = T16709[6'h27:6'h27];
  assign T16713 = T10817[1'h0:1'h0];
  assign T16714 = T10817[1'h1:1'h1];
  assign T16715 = T10817[2'h2:2'h2];
  assign T16716 = T10817[2'h3:2'h3];
  assign T16717 = T10817[3'h4:3'h4];
  assign T16718 = T10817[3'h5:3'h5];
  assign T16719 = T10817[3'h6:3'h6];
  assign T16720 = T15743[6'h2e:6'h2e];
  assign T16721 = T10817[3'h7:3'h7];
  assign T16722 = T18696 ? T17717 : T16723;
  assign T16723 = T17716 ? T17288 : T16724;
  assign T16724 = T17287 ? T17021 : T16725;
  assign T16725 = T17020 ? T16876 : T16726;
  assign T16726 = T16875 ? T16803 : T16727;
  assign T16727 = T16802 ? T16766 : T16728;
  assign T16728 = T16765 ? T16747 : T16729;
  assign T16729 = T16746 ? T16737 : twiddle4_2_256_real;
  assign twiddle4_2_256_real = T16732 + T16730;
  assign T16730 = $signed(T16731) / $signed(22'h100000);
  assign T16731 = $signed(32'h40000000) * $signed(16'h0);
  assign T16732 = {T16735, T16733};
  assign T16733 = $signed(T16734) / $signed(22'h100000);
  assign T16734 = $signed(1'h0) * $signed(16'h1);
  assign T16735 = T16736 ? 31'h7fffffff : 31'h0;
  assign T16736 = T16733[5'h10:5'h10];
  assign T16737 = {T16745, twiddle4_2_257_real};
  assign twiddle4_2_257_real = T16740 + T16738;
  assign T16738 = $signed(T16739) / $signed(22'h100000);
  assign T16739 = $signed(31'h3fffb10b) * $signed(16'h0);
  assign T16740 = {T16743, T16741};
  assign T16741 = $signed(T16742) / $signed(22'h100000);
  assign T16742 = $signed(24'h9b783d) * $signed(16'h1);
  assign T16743 = T16744 ? 7'h7f : 7'h0;
  assign T16744 = T16741[6'h27:6'h27];
  assign T16745 = twiddle4_2_257_real[6'h2e:6'h2e];
  assign T16746 = T10817[1'h0:1'h0];
  assign T16747 = {T16764, T16748};
  assign T16748 = T16763 ? twiddle4_2_259_real : twiddle4_2_258_real;
  assign twiddle4_2_258_real = T16751 + T16749;
  assign T16749 = $signed(T16750) / $signed(22'h100000);
  assign T16750 = $signed(31'h3ffec42d) * $signed(16'h0);
  assign T16751 = {T16754, T16752};
  assign T16752 = $signed(T16753) / $signed(22'h100000);
  assign T16753 = $signed(25'h136f171) * $signed(16'h1);
  assign T16754 = T16755 ? 6'h3f : 6'h0;
  assign T16755 = T16752[6'h28:6'h28];
  assign twiddle4_2_259_real = T16758 + T16756;
  assign T16756 = $signed(T16757) / $signed(22'h100000);
  assign T16757 = $signed(31'h3ffd3968) * $signed(16'h0);
  assign T16758 = {T16761, T16759};
  assign T16759 = $signed(T16760) / $signed(22'h100000);
  assign T16760 = $signed(26'h2d26c95) * $signed(16'h1);
  assign T16761 = T16762 ? 5'h1f : 5'h0;
  assign T16762 = T16759[6'h29:6'h29];
  assign T16763 = T10817[1'h0:1'h0];
  assign T16764 = T16748[6'h2e:6'h2e];
  assign T16765 = T10817[1'h1:1'h1];
  assign T16766 = {T16801, T16767};
  assign T16767 = T16800 ? T16784 : T16768;
  assign T16768 = T16783 ? twiddle4_2_261_real : twiddle4_2_260_real;
  assign twiddle4_2_260_real = T16771 + T16769;
  assign T16769 = $signed(T16770) / $signed(22'h100000);
  assign T16770 = $signed(31'h3ffb10c1) * $signed(16'h0);
  assign T16771 = {T16774, T16772};
  assign T16772 = $signed(T16773) / $signed(22'h100000);
  assign T16773 = $signed(26'h26deaa1) * $signed(16'h1);
  assign T16774 = T16775 ? 5'h1f : 5'h0;
  assign T16775 = T16772[6'h29:6'h29];
  assign twiddle4_2_261_real = T16778 + T16776;
  assign T16776 = $signed(T16777) / $signed(22'h100000);
  assign T16777 = $signed(31'h3ff84a3b) * $signed(16'h0);
  assign T16778 = {T16781, T16779};
  assign T16779 = $signed(T16780) / $signed(22'h100000);
  assign T16780 = $signed(26'h2096c8d) * $signed(16'h1);
  assign T16781 = T16782 ? 5'h1f : 5'h0;
  assign T16782 = T16779[6'h29:6'h29];
  assign T16783 = T10817[1'h0:1'h0];
  assign T16784 = T16799 ? twiddle4_2_263_real : twiddle4_2_262_real;
  assign twiddle4_2_262_real = T16787 + T16785;
  assign T16785 = $signed(T16786) / $signed(22'h100000);
  assign T16786 = $signed(31'h3ff4e5df) * $signed(16'h0);
  assign T16787 = {T16790, T16788};
  assign T16788 = $signed(T16789) / $signed(22'h100000);
  assign T16789 = $signed(27'h5a4f352) * $signed(16'h1);
  assign T16790 = T16791 ? 4'hf : 4'h0;
  assign T16791 = T16788[6'h2a:6'h2a];
  assign twiddle4_2_263_real = T16794 + T16792;
  assign T16792 = $signed(T16793) / $signed(22'h100000);
  assign T16793 = $signed(31'h3ff0e3b5) * $signed(16'h0);
  assign T16794 = {T16797, T16795};
  assign T16795 = $signed(T16796) / $signed(22'h100000);
  assign T16796 = $signed(27'h5407fe6) * $signed(16'h1);
  assign T16797 = T16798 ? 4'hf : 4'h0;
  assign T16798 = T16795[6'h2a:6'h2a];
  assign T16799 = T10817[1'h0:1'h0];
  assign T16800 = T10817[1'h1:1'h1];
  assign T16801 = T16767[6'h2e:6'h2e];
  assign T16802 = T10817[2'h2:2'h2];
  assign T16803 = {T16874, T16804};
  assign T16804 = T16873 ? T16839 : T16805;
  assign T16805 = T16838 ? T16822 : T16806;
  assign T16806 = T16821 ? twiddle4_2_265_real : twiddle4_2_264_real;
  assign twiddle4_2_264_real = T16809 + T16807;
  assign T16807 = $signed(T16808) / $signed(22'h100000);
  assign T16808 = $signed(31'h3fec43c6) * $signed(16'h0);
  assign T16809 = {T16812, T16810};
  assign T16810 = $signed(T16811) / $signed(22'h100000);
  assign T16811 = $signed(27'h4dc1342) * $signed(16'h1);
  assign T16812 = T16813 ? 4'hf : 4'h0;
  assign T16813 = T16810[6'h2a:6'h2a];
  assign twiddle4_2_265_real = T16816 + T16814;
  assign T16814 = $signed(T16815) / $signed(22'h100000);
  assign T16815 = $signed(31'h3fe7061f) * $signed(16'h0);
  assign T16816 = {T16819, T16817};
  assign T16817 = $signed(T16818) / $signed(22'h100000);
  assign T16818 = $signed(27'h477ae5e) * $signed(16'h1);
  assign T16819 = T16820 ? 4'hf : 4'h0;
  assign T16820 = T16817[6'h2a:6'h2a];
  assign T16821 = T10817[1'h0:1'h0];
  assign T16822 = T16837 ? twiddle4_2_267_real : twiddle4_2_266_real;
  assign twiddle4_2_266_real = T16825 + T16823;
  assign T16823 = $signed(T16824) / $signed(22'h100000);
  assign T16824 = $signed(31'h3fe12acb) * $signed(16'h0);
  assign T16825 = {T16828, T16826};
  assign T16826 = $signed(T16827) / $signed(22'h100000);
  assign T16827 = $signed(27'h4135231) * $signed(16'h1);
  assign T16828 = T16829 ? 4'hf : 4'h0;
  assign T16829 = T16826[6'h2a:6'h2a];
  assign twiddle4_2_267_real = T16832 + T16830;
  assign T16830 = $signed(T16831) / $signed(22'h100000);
  assign T16831 = $signed(31'h3fdab1d9) * $signed(16'h0);
  assign T16832 = {T16835, T16833};
  assign T16833 = $signed(T16834) / $signed(22'h100000);
  assign T16834 = $signed(28'hbaeffb3) * $signed(16'h1);
  assign T16835 = T16836 ? 3'h7 : 3'h0;
  assign T16836 = T16833[6'h2b:6'h2b];
  assign T16837 = T10817[1'h0:1'h0];
  assign T16838 = T10817[1'h1:1'h1];
  assign T16839 = T16872 ? T16856 : T16840;
  assign T16840 = T16855 ? twiddle4_2_269_real : twiddle4_2_268_real;
  assign twiddle4_2_268_real = T16843 + T16841;
  assign T16841 = $signed(T16842) / $signed(22'h100000);
  assign T16842 = $signed(31'h3fd39b5a) * $signed(16'h0);
  assign T16843 = {T16846, T16844};
  assign T16844 = $signed(T16845) / $signed(22'h100000);
  assign T16845 = $signed(28'hb4ab7dc) * $signed(16'h1);
  assign T16846 = T16847 ? 3'h7 : 3'h0;
  assign T16847 = T16844[6'h2b:6'h2b];
  assign twiddle4_2_269_real = T16850 + T16848;
  assign T16848 = $signed(T16849) / $signed(22'h100000);
  assign T16849 = $signed(31'h3fcbe75e) * $signed(16'h0);
  assign T16850 = {T16853, T16851};
  assign T16851 = $signed(T16852) / $signed(22'h100000);
  assign T16852 = $signed(28'hae67ba2) * $signed(16'h1);
  assign T16853 = T16854 ? 3'h7 : 3'h0;
  assign T16854 = T16851[6'h2b:6'h2b];
  assign T16855 = T10817[1'h0:1'h0];
  assign T16856 = T16871 ? twiddle4_2_271_real : twiddle4_2_270_real;
  assign twiddle4_2_270_real = T16859 + T16857;
  assign T16857 = $signed(T16858) / $signed(22'h100000);
  assign T16858 = $signed(31'h3fc395f9) * $signed(16'h0);
  assign T16859 = {T16862, T16860};
  assign T16860 = $signed(T16861) / $signed(22'h100000);
  assign T16861 = $signed(28'ha824bfe) * $signed(16'h1);
  assign T16862 = T16863 ? 3'h7 : 3'h0;
  assign T16863 = T16860[6'h2b:6'h2b];
  assign twiddle4_2_271_real = T16866 + T16864;
  assign T16864 = $signed(T16865) / $signed(22'h100000);
  assign T16865 = $signed(31'h3fbaa73f) * $signed(16'h0);
  assign T16866 = {T16869, T16867};
  assign T16867 = $signed(T16868) / $signed(22'h100000);
  assign T16868 = $signed(28'ha1e29e6) * $signed(16'h1);
  assign T16869 = T16870 ? 3'h7 : 3'h0;
  assign T16870 = T16867[6'h2b:6'h2b];
  assign T16871 = T10817[1'h0:1'h0];
  assign T16872 = T10817[1'h1:1'h1];
  assign T16873 = T10817[2'h2:2'h2];
  assign T16874 = T16804[6'h2e:6'h2e];
  assign T16875 = T10817[2'h3:2'h3];
  assign T16876 = {T17019, T16877};
  assign T16877 = T17018 ? T16948 : T16878;
  assign T16878 = T16947 ? T16913 : T16879;
  assign T16879 = T16912 ? T16896 : T16880;
  assign T16880 = T16895 ? twiddle4_2_273_real : twiddle4_2_272_real;
  assign twiddle4_2_272_real = T16883 + T16881;
  assign T16881 = $signed(T16882) / $signed(22'h100000);
  assign T16882 = $signed(31'h3fb11b47) * $signed(16'h0);
  assign T16883 = {T16886, T16884};
  assign T16884 = $signed(T16885) / $signed(22'h100000);
  assign T16885 = $signed(28'h9ba1651) * $signed(16'h1);
  assign T16886 = T16887 ? 3'h7 : 3'h0;
  assign T16887 = T16884[6'h2b:6'h2b];
  assign twiddle4_2_273_real = T16890 + T16888;
  assign T16888 = $signed(T16889) / $signed(22'h100000);
  assign T16889 = $signed(31'h3fa6f228) * $signed(16'h0);
  assign T16890 = {T16893, T16891};
  assign T16891 = $signed(T16892) / $signed(22'h100000);
  assign T16892 = $signed(28'h9561237) * $signed(16'h1);
  assign T16893 = T16894 ? 3'h7 : 3'h0;
  assign T16894 = T16891[6'h2b:6'h2b];
  assign T16895 = T10817[1'h0:1'h0];
  assign T16896 = T16911 ? twiddle4_2_275_real : twiddle4_2_274_real;
  assign twiddle4_2_274_real = T16899 + T16897;
  assign T16897 = $signed(T16898) / $signed(22'h100000);
  assign T16898 = $signed(31'h3f9c2bfa) * $signed(16'h0);
  assign T16899 = {T16902, T16900};
  assign T16900 = $signed(T16901) / $signed(22'h100000);
  assign T16901 = $signed(28'h8f21e8f) * $signed(16'h1);
  assign T16902 = T16903 ? 3'h7 : 3'h0;
  assign T16903 = T16900[6'h2b:6'h2b];
  assign twiddle4_2_275_real = T16906 + T16904;
  assign T16904 = $signed(T16905) / $signed(22'h100000);
  assign T16905 = $signed(31'h3f90c8d9) * $signed(16'h0);
  assign T16906 = {T16909, T16907};
  assign T16907 = $signed(T16908) / $signed(22'h100000);
  assign T16908 = $signed(28'h88e3c4e) * $signed(16'h1);
  assign T16909 = T16910 ? 3'h7 : 3'h0;
  assign T16910 = T16907[6'h2b:6'h2b];
  assign T16911 = T10817[1'h0:1'h0];
  assign T16912 = T10817[1'h1:1'h1];
  assign T16913 = T16946 ? T16930 : T16914;
  assign T16914 = T16929 ? twiddle4_2_277_real : twiddle4_2_276_real;
  assign twiddle4_2_276_real = T16917 + T16915;
  assign T16915 = $signed(T16916) / $signed(22'h100000);
  assign T16916 = $signed(31'h3f84c8e1) * $signed(16'h0);
  assign T16917 = {T16920, T16918};
  assign T16918 = $signed(T16919) / $signed(22'h100000);
  assign T16919 = $signed(28'h82a6c6b) * $signed(16'h1);
  assign T16920 = T16921 ? 3'h7 : 3'h0;
  assign T16921 = T16918[6'h2b:6'h2b];
  assign twiddle4_2_277_real = T16924 + T16922;
  assign T16922 = $signed(T16923) / $signed(22'h100000);
  assign T16923 = $signed(31'h3f782c2f) * $signed(16'h0);
  assign T16924 = {T16927, T16925};
  assign T16925 = $signed(T16926) / $signed(22'h100000);
  assign T16926 = $signed(29'h17c6afdd) * $signed(16'h1);
  assign T16927 = T16928 ? 2'h3 : 2'h0;
  assign T16928 = T16925[6'h2c:6'h2c];
  assign T16929 = T10817[1'h0:1'h0];
  assign T16930 = T16945 ? twiddle4_2_279_real : twiddle4_2_278_real;
  assign twiddle4_2_278_real = T16933 + T16931;
  assign T16931 = $signed(T16932) / $signed(22'h100000);
  assign T16932 = $signed(31'h3f6af2e3) * $signed(16'h0);
  assign T16933 = {T16936, T16934};
  assign T16934 = $signed(T16935) / $signed(22'h100000);
  assign T16935 = $signed(29'h17630799) * $signed(16'h1);
  assign T16936 = T16937 ? 2'h3 : 2'h0;
  assign T16937 = T16934[6'h2c:6'h2c];
  assign twiddle4_2_279_real = T16940 + T16938;
  assign T16938 = $signed(T16939) / $signed(22'h100000);
  assign T16939 = $signed(31'h3f5d1d1c) * $signed(16'h0);
  assign T16940 = {T16943, T16941};
  assign T16941 = $signed(T16942) / $signed(22'h100000);
  assign T16942 = $signed(29'h16ff7496) * $signed(16'h1);
  assign T16943 = T16944 ? 2'h3 : 2'h0;
  assign T16944 = T16941[6'h2c:6'h2c];
  assign T16945 = T10817[1'h0:1'h0];
  assign T16946 = T10817[1'h1:1'h1];
  assign T16947 = T10817[2'h2:2'h2];
  assign T16948 = T17017 ? T16983 : T16949;
  assign T16949 = T16982 ? T16966 : T16950;
  assign T16950 = T16965 ? twiddle4_2_281_real : twiddle4_2_280_real;
  assign twiddle4_2_280_real = T16953 + T16951;
  assign T16951 = $signed(T16952) / $signed(22'h100000);
  assign T16952 = $signed(31'h3f4eaafe) * $signed(16'h0);
  assign T16953 = {T16956, T16954};
  assign T16954 = $signed(T16955) / $signed(22'h100000);
  assign T16955 = $signed(29'h169bf7c9) * $signed(16'h1);
  assign T16956 = T16957 ? 2'h3 : 2'h0;
  assign T16957 = T16954[6'h2c:6'h2c];
  assign twiddle4_2_281_real = T16960 + T16958;
  assign T16958 = $signed(T16959) / $signed(22'h100000);
  assign T16959 = $signed(31'h3f3f9cab) * $signed(16'h0);
  assign T16960 = {T16963, T16961};
  assign T16961 = $signed(T16962) / $signed(22'h100000);
  assign T16962 = $signed(29'h16389228) * $signed(16'h1);
  assign T16963 = T16964 ? 2'h3 : 2'h0;
  assign T16964 = T16961[6'h2c:6'h2c];
  assign T16965 = T10817[1'h0:1'h0];
  assign T16966 = T16981 ? twiddle4_2_283_real : twiddle4_2_282_real;
  assign twiddle4_2_282_real = T16969 + T16967;
  assign T16967 = $signed(T16968) / $signed(22'h100000);
  assign T16968 = $signed(31'h3f2ff249) * $signed(16'h0);
  assign T16969 = {T16972, T16970};
  assign T16970 = $signed(T16971) / $signed(22'h100000);
  assign T16971 = $signed(29'h15d544a8) * $signed(16'h1);
  assign T16972 = T16973 ? 2'h3 : 2'h0;
  assign T16973 = T16970[6'h2c:6'h2c];
  assign twiddle4_2_283_real = T16976 + T16974;
  assign T16974 = $signed(T16975) / $signed(22'h100000);
  assign T16975 = $signed(31'h3f1fabff) * $signed(16'h0);
  assign T16976 = {T16979, T16977};
  assign T16977 = $signed(T16978) / $signed(22'h100000);
  assign T16978 = $signed(29'h1572103e) * $signed(16'h1);
  assign T16979 = T16980 ? 2'h3 : 2'h0;
  assign T16980 = T16977[6'h2c:6'h2c];
  assign T16981 = T10817[1'h0:1'h0];
  assign T16982 = T10817[1'h1:1'h1];
  assign T16983 = T17016 ? T17000 : T16984;
  assign T16984 = T16999 ? twiddle4_2_285_real : twiddle4_2_284_real;
  assign twiddle4_2_284_real = T16987 + T16985;
  assign T16985 = $signed(T16986) / $signed(22'h100000);
  assign T16986 = $signed(31'h3f0ec9f4) * $signed(16'h0);
  assign T16987 = {T16990, T16988};
  assign T16988 = $signed(T16989) / $signed(22'h100000);
  assign T16989 = $signed(29'h150ef5de) * $signed(16'h1);
  assign T16990 = T16991 ? 2'h3 : 2'h0;
  assign T16991 = T16988[6'h2c:6'h2c];
  assign twiddle4_2_285_real = T16994 + T16992;
  assign T16992 = $signed(T16993) / $signed(22'h100000);
  assign T16993 = $signed(31'h3efd4c53) * $signed(16'h0);
  assign T16994 = {T16997, T16995};
  assign T16995 = $signed(T16996) / $signed(22'h100000);
  assign T16996 = $signed(29'h14abf67e) * $signed(16'h1);
  assign T16997 = T16998 ? 2'h3 : 2'h0;
  assign T16998 = T16995[6'h2c:6'h2c];
  assign T16999 = T10817[1'h0:1'h0];
  assign T17000 = T17015 ? twiddle4_2_287_real : twiddle4_2_286_real;
  assign twiddle4_2_286_real = T17003 + T17001;
  assign T17001 = $signed(T17002) / $signed(22'h100000);
  assign T17002 = $signed(31'h3eeb3347) * $signed(16'h0);
  assign T17003 = {T17006, T17004};
  assign T17004 = $signed(T17005) / $signed(22'h100000);
  assign T17005 = $signed(29'h14491311) * $signed(16'h1);
  assign T17006 = T17007 ? 2'h3 : 2'h0;
  assign T17007 = T17004[6'h2c:6'h2c];
  assign twiddle4_2_287_real = T17010 + T17008;
  assign T17008 = $signed(T17009) / $signed(22'h100000);
  assign T17009 = $signed(31'h3ed87efb) * $signed(16'h0);
  assign T17010 = {T17013, T17011};
  assign T17011 = $signed(T17012) / $signed(22'h100000);
  assign T17012 = $signed(29'h13e64c8c) * $signed(16'h1);
  assign T17013 = T17014 ? 2'h3 : 2'h0;
  assign T17014 = T17011[6'h2c:6'h2c];
  assign T17015 = T10817[1'h0:1'h0];
  assign T17016 = T10817[1'h1:1'h1];
  assign T17017 = T10817[2'h2:2'h2];
  assign T17018 = T10817[2'h3:2'h3];
  assign T17019 = T16877[6'h2e:6'h2e];
  assign T17020 = T10817[3'h4:3'h4];
  assign T17021 = {T17286, T17022};
  assign T17022 = T17285 ? T17159 : T17023;
  assign T17023 = T17158 ? T17094 : T17024;
  assign T17024 = T17093 ? T17059 : T17025;
  assign T17025 = T17058 ? T17042 : T17026;
  assign T17026 = T17041 ? twiddle4_2_289_real : twiddle4_2_288_real;
  assign twiddle4_2_288_real = T17029 + T17027;
  assign T17027 = $signed(T17028) / $signed(22'h100000);
  assign T17028 = $signed(31'h3ec52f9f) * $signed(16'h0);
  assign T17029 = {T17032, T17030};
  assign T17030 = $signed(T17031) / $signed(22'h100000);
  assign T17031 = $signed(29'h1383a3e2) * $signed(16'h1);
  assign T17032 = T17033 ? 2'h3 : 2'h0;
  assign T17033 = T17030[6'h2c:6'h2c];
  assign twiddle4_2_289_real = T17036 + T17034;
  assign T17034 = $signed(T17035) / $signed(22'h100000);
  assign T17035 = $signed(31'h3eb14562) * $signed(16'h0);
  assign T17036 = {T17039, T17037};
  assign T17037 = $signed(T17038) / $signed(22'h100000);
  assign T17038 = $signed(29'h13211a07) * $signed(16'h1);
  assign T17039 = T17040 ? 2'h3 : 2'h0;
  assign T17040 = T17037[6'h2c:6'h2c];
  assign T17041 = T10817[1'h0:1'h0];
  assign T17042 = T17057 ? twiddle4_2_291_real : twiddle4_2_290_real;
  assign twiddle4_2_290_real = T17045 + T17043;
  assign T17043 = $signed(T17044) / $signed(22'h100000);
  assign T17044 = $signed(31'h3e9cc076) * $signed(16'h0);
  assign T17045 = {T17048, T17046};
  assign T17046 = $signed(T17047) / $signed(22'h100000);
  assign T17047 = $signed(29'h12beafee) * $signed(16'h1);
  assign T17048 = T17049 ? 2'h3 : 2'h0;
  assign T17049 = T17046[6'h2c:6'h2c];
  assign twiddle4_2_291_real = T17052 + T17050;
  assign T17050 = $signed(T17051) / $signed(22'h100000);
  assign T17051 = $signed(31'h3e87a10b) * $signed(16'h0);
  assign T17052 = {T17055, T17053};
  assign T17053 = $signed(T17054) / $signed(22'h100000);
  assign T17054 = $signed(29'h125c6689) * $signed(16'h1);
  assign T17055 = T17056 ? 2'h3 : 2'h0;
  assign T17056 = T17053[6'h2c:6'h2c];
  assign T17057 = T10817[1'h0:1'h0];
  assign T17058 = T10817[1'h1:1'h1];
  assign T17059 = T17092 ? T17076 : T17060;
  assign T17060 = T17075 ? twiddle4_2_293_real : twiddle4_2_292_real;
  assign twiddle4_2_292_real = T17063 + T17061;
  assign T17061 = $signed(T17062) / $signed(22'h100000);
  assign T17062 = $signed(31'h3e71e758) * $signed(16'h0);
  assign T17063 = {T17066, T17064};
  assign T17064 = $signed(T17065) / $signed(22'h100000);
  assign T17065 = $signed(29'h11fa3ecb) * $signed(16'h1);
  assign T17066 = T17067 ? 2'h3 : 2'h0;
  assign T17067 = T17064[6'h2c:6'h2c];
  assign twiddle4_2_293_real = T17070 + T17068;
  assign T17068 = $signed(T17069) / $signed(22'h100000);
  assign T17069 = $signed(31'h3e5b9392) * $signed(16'h0);
  assign T17070 = {T17073, T17071};
  assign T17071 = $signed(T17072) / $signed(22'h100000);
  assign T17072 = $signed(29'h119839a7) * $signed(16'h1);
  assign T17073 = T17074 ? 2'h3 : 2'h0;
  assign T17074 = T17071[6'h2c:6'h2c];
  assign T17075 = T10817[1'h0:1'h0];
  assign T17076 = T17091 ? twiddle4_2_295_real : twiddle4_2_294_real;
  assign twiddle4_2_294_real = T17079 + T17077;
  assign T17077 = $signed(T17078) / $signed(22'h100000);
  assign T17078 = $signed(31'h3e44a5ee) * $signed(16'h0);
  assign T17079 = {T17082, T17080};
  assign T17080 = $signed(T17081) / $signed(22'h100000);
  assign T17081 = $signed(29'h1136580e) * $signed(16'h1);
  assign T17082 = T17083 ? 2'h3 : 2'h0;
  assign T17083 = T17080[6'h2c:6'h2c];
  assign twiddle4_2_295_real = T17086 + T17084;
  assign T17084 = $signed(T17085) / $signed(22'h100000);
  assign T17085 = $signed(31'h3e2d1ea7) * $signed(16'h0);
  assign T17086 = {T17089, T17087};
  assign T17087 = $signed(T17088) / $signed(22'h100000);
  assign T17088 = $signed(29'h10d49af1) * $signed(16'h1);
  assign T17089 = T17090 ? 2'h3 : 2'h0;
  assign T17090 = T17087[6'h2c:6'h2c];
  assign T17091 = T10817[1'h0:1'h0];
  assign T17092 = T10817[1'h1:1'h1];
  assign T17093 = T10817[2'h2:2'h2];
  assign T17094 = T17157 ? T17127 : T17095;
  assign T17095 = T17126 ? T17112 : T17096;
  assign T17096 = T17111 ? twiddle4_2_297_real : twiddle4_2_296_real;
  assign twiddle4_2_296_real = T17099 + T17097;
  assign T17097 = $signed(T17098) / $signed(22'h100000);
  assign T17098 = $signed(31'h3e14fdf7) * $signed(16'h0);
  assign T17099 = {T17102, T17100};
  assign T17100 = $signed(T17101) / $signed(22'h100000);
  assign T17101 = $signed(29'h10730343) * $signed(16'h1);
  assign T17102 = T17103 ? 2'h3 : 2'h0;
  assign T17103 = T17100[6'h2c:6'h2c];
  assign twiddle4_2_297_real = T17106 + T17104;
  assign T17104 = $signed(T17105) / $signed(22'h100000);
  assign T17105 = $signed(31'h3dfc4418) * $signed(16'h0);
  assign T17106 = {T17109, T17107};
  assign T17107 = $signed(T17108) / $signed(22'h100000);
  assign T17108 = $signed(29'h101191f3) * $signed(16'h1);
  assign T17109 = T17110 ? 2'h3 : 2'h0;
  assign T17110 = T17107[6'h2c:6'h2c];
  assign T17111 = T10817[1'h0:1'h0];
  assign T17112 = T17125 ? twiddle4_2_299_real : twiddle4_2_298_real;
  assign twiddle4_2_298_real = T17115 + T17113;
  assign T17113 = $signed(T17114) / $signed(22'h100000);
  assign T17114 = $signed(31'h3de2f147) * $signed(16'h0);
  assign T17115 = {T17118, T17116};
  assign T17116 = $signed(T17117) / $signed(22'h100000);
  assign T17117 = $signed(30'h2fb047f2) * $signed(16'h1);
  assign T17118 = T17116[6'h2d:6'h2d];
  assign twiddle4_2_299_real = T17121 + T17119;
  assign T17119 = $signed(T17120) / $signed(22'h100000);
  assign T17120 = $signed(31'h3dc905c4) * $signed(16'h0);
  assign T17121 = {T17124, T17122};
  assign T17122 = $signed(T17123) / $signed(22'h100000);
  assign T17123 = $signed(30'h2f4f2631) * $signed(16'h1);
  assign T17124 = T17122[6'h2d:6'h2d];
  assign T17125 = T10817[1'h0:1'h0];
  assign T17126 = T10817[1'h1:1'h1];
  assign T17127 = T17156 ? T17142 : T17128;
  assign T17128 = T17141 ? twiddle4_2_301_real : twiddle4_2_300_real;
  assign twiddle4_2_300_real = T17131 + T17129;
  assign T17129 = $signed(T17130) / $signed(22'h100000);
  assign T17130 = $signed(31'h3dae81ce) * $signed(16'h0);
  assign T17131 = {T17134, T17132};
  assign T17132 = $signed(T17133) / $signed(22'h100000);
  assign T17133 = $signed(30'h2eee2d9e) * $signed(16'h1);
  assign T17134 = T17132[6'h2d:6'h2d];
  assign twiddle4_2_301_real = T17137 + T17135;
  assign T17135 = $signed(T17136) / $signed(22'h100000);
  assign T17136 = $signed(31'h3d9365a7) * $signed(16'h0);
  assign T17137 = {T17140, T17138};
  assign T17138 = $signed(T17139) / $signed(22'h100000);
  assign T17139 = $signed(30'h2e8d5f29) * $signed(16'h1);
  assign T17140 = T17138[6'h2d:6'h2d];
  assign T17141 = T10817[1'h0:1'h0];
  assign T17142 = T17155 ? twiddle4_2_303_real : twiddle4_2_302_real;
  assign twiddle4_2_302_real = T17145 + T17143;
  assign T17143 = $signed(T17144) / $signed(22'h100000);
  assign T17144 = $signed(31'h3d77b191) * $signed(16'h0);
  assign T17145 = {T17148, T17146};
  assign T17146 = $signed(T17147) / $signed(22'h100000);
  assign T17147 = $signed(30'h2e2cbbc1) * $signed(16'h1);
  assign T17148 = T17146[6'h2d:6'h2d];
  assign twiddle4_2_303_real = T17151 + T17149;
  assign T17149 = $signed(T17150) / $signed(22'h100000);
  assign T17150 = $signed(31'h3d5b65d1) * $signed(16'h0);
  assign T17151 = {T17154, T17152};
  assign T17152 = $signed(T17153) / $signed(22'h100000);
  assign T17153 = $signed(30'h2dcc4455) * $signed(16'h1);
  assign T17154 = T17152[6'h2d:6'h2d];
  assign T17155 = T10817[1'h0:1'h0];
  assign T17156 = T10817[1'h1:1'h1];
  assign T17157 = T10817[2'h2:2'h2];
  assign T17158 = T10817[2'h3:2'h3];
  assign T17159 = T17284 ? T17222 : T17160;
  assign T17160 = T17221 ? T17191 : T17161;
  assign T17161 = T17190 ? T17176 : T17162;
  assign T17162 = T17175 ? twiddle4_2_305_real : twiddle4_2_304_real;
  assign twiddle4_2_304_real = T17165 + T17163;
  assign T17163 = $signed(T17164) / $signed(22'h100000);
  assign T17164 = $signed(31'h3d3e82ad) * $signed(16'h0);
  assign T17165 = {T17168, T17166};
  assign T17166 = $signed(T17167) / $signed(22'h100000);
  assign T17167 = $signed(30'h2d6bf9d2) * $signed(16'h1);
  assign T17168 = T17166[6'h2d:6'h2d];
  assign twiddle4_2_305_real = T17171 + T17169;
  assign T17169 = $signed(T17170) / $signed(22'h100000);
  assign T17170 = $signed(31'h3d21086c) * $signed(16'h0);
  assign T17171 = {T17174, T17172};
  assign T17172 = $signed(T17173) / $signed(22'h100000);
  assign T17173 = $signed(30'h2d0bdd26) * $signed(16'h1);
  assign T17174 = T17172[6'h2d:6'h2d];
  assign T17175 = T10817[1'h0:1'h0];
  assign T17176 = T17189 ? twiddle4_2_307_real : twiddle4_2_306_real;
  assign twiddle4_2_306_real = T17179 + T17177;
  assign T17177 = $signed(T17178) / $signed(22'h100000);
  assign T17178 = $signed(31'h3d02f756) * $signed(16'h0);
  assign T17179 = {T17182, T17180};
  assign T17180 = $signed(T17181) / $signed(22'h100000);
  assign T17181 = $signed(30'h2cabef3e) * $signed(16'h1);
  assign T17182 = T17180[6'h2d:6'h2d];
  assign twiddle4_2_307_real = T17185 + T17183;
  assign T17183 = $signed(T17184) / $signed(22'h100000);
  assign T17184 = $signed(31'h3ce44fb6) * $signed(16'h0);
  assign T17185 = {T17188, T17186};
  assign T17186 = $signed(T17187) / $signed(22'h100000);
  assign T17187 = $signed(30'h2c4c3106) * $signed(16'h1);
  assign T17188 = T17186[6'h2d:6'h2d];
  assign T17189 = T10817[1'h0:1'h0];
  assign T17190 = T10817[1'h1:1'h1];
  assign T17191 = T17220 ? T17206 : T17192;
  assign T17192 = T17205 ? twiddle4_2_309_real : twiddle4_2_308_real;
  assign twiddle4_2_308_real = T17195 + T17193;
  assign T17193 = $signed(T17194) / $signed(22'h100000);
  assign T17194 = $signed(31'h3cc511d8) * $signed(16'h0);
  assign T17195 = {T17198, T17196};
  assign T17196 = $signed(T17197) / $signed(22'h100000);
  assign T17197 = $signed(30'h2beca36c) * $signed(16'h1);
  assign T17198 = T17196[6'h2d:6'h2d];
  assign twiddle4_2_309_real = T17201 + T17199;
  assign T17199 = $signed(T17200) / $signed(22'h100000);
  assign T17200 = $signed(31'h3ca53e08) * $signed(16'h0);
  assign T17201 = {T17204, T17202};
  assign T17202 = $signed(T17203) / $signed(22'h100000);
  assign T17203 = $signed(30'h2b8d475b) * $signed(16'h1);
  assign T17204 = T17202[6'h2d:6'h2d];
  assign T17205 = T10817[1'h0:1'h0];
  assign T17206 = T17219 ? twiddle4_2_311_real : twiddle4_2_310_real;
  assign twiddle4_2_310_real = T17209 + T17207;
  assign T17207 = $signed(T17208) / $signed(22'h100000);
  assign T17208 = $signed(31'h3c84d496) * $signed(16'h0);
  assign T17209 = {T17212, T17210};
  assign T17210 = $signed(T17211) / $signed(22'h100000);
  assign T17211 = $signed(30'h2b2e1dbe) * $signed(16'h1);
  assign T17212 = T17210[6'h2d:6'h2d];
  assign twiddle4_2_311_real = T17215 + T17213;
  assign T17213 = $signed(T17214) / $signed(22'h100000);
  assign T17214 = $signed(31'h3c63d5d0) * $signed(16'h0);
  assign T17215 = {T17218, T17216};
  assign T17216 = $signed(T17217) / $signed(22'h100000);
  assign T17217 = $signed(30'h2acf2780) * $signed(16'h1);
  assign T17218 = T17216[6'h2d:6'h2d];
  assign T17219 = T10817[1'h0:1'h0];
  assign T17220 = T10817[1'h1:1'h1];
  assign T17221 = T10817[2'h2:2'h2];
  assign T17222 = T17283 ? T17253 : T17223;
  assign T17223 = T17252 ? T17238 : T17224;
  assign T17224 = T17237 ? twiddle4_2_313_real : twiddle4_2_312_real;
  assign twiddle4_2_312_real = T17227 + T17225;
  assign T17225 = $signed(T17226) / $signed(22'h100000);
  assign T17226 = $signed(31'h3c424209) * $signed(16'h0);
  assign T17227 = {T17230, T17228};
  assign T17228 = $signed(T17229) / $signed(22'h100000);
  assign T17229 = $signed(30'h2a70658b) * $signed(16'h1);
  assign T17230 = T17228[6'h2d:6'h2d];
  assign twiddle4_2_313_real = T17233 + T17231;
  assign T17231 = $signed(T17232) / $signed(22'h100000);
  assign T17232 = $signed(31'h3c201994) * $signed(16'h0);
  assign T17233 = {T17236, T17234};
  assign T17234 = $signed(T17235) / $signed(22'h100000);
  assign T17235 = $signed(30'h2a11d8c9) * $signed(16'h1);
  assign T17236 = T17234[6'h2d:6'h2d];
  assign T17237 = T10817[1'h0:1'h0];
  assign T17238 = T17251 ? twiddle4_2_315_real : twiddle4_2_314_real;
  assign twiddle4_2_314_real = T17241 + T17239;
  assign T17239 = $signed(T17240) / $signed(22'h100000);
  assign T17240 = $signed(31'h3bfd5cc4) * $signed(16'h0);
  assign T17241 = {T17244, T17242};
  assign T17242 = $signed(T17243) / $signed(22'h100000);
  assign T17243 = $signed(30'h29b38223) * $signed(16'h1);
  assign T17244 = T17242[6'h2d:6'h2d];
  assign twiddle4_2_315_real = T17247 + T17245;
  assign T17245 = $signed(T17246) / $signed(22'h100000);
  assign T17246 = $signed(31'h3bda0bef) * $signed(16'h0);
  assign T17247 = {T17250, T17248};
  assign T17248 = $signed(T17249) / $signed(22'h100000);
  assign T17249 = $signed(30'h29556283) * $signed(16'h1);
  assign T17250 = T17248[6'h2d:6'h2d];
  assign T17251 = T10817[1'h0:1'h0];
  assign T17252 = T10817[1'h1:1'h1];
  assign T17253 = T17282 ? T17268 : T17254;
  assign T17254 = T17267 ? twiddle4_2_317_real : twiddle4_2_316_real;
  assign twiddle4_2_316_real = T17257 + T17255;
  assign T17255 = $signed(T17256) / $signed(22'h100000);
  assign T17256 = $signed(31'h3bb6276d) * $signed(16'h0);
  assign T17257 = {T17260, T17258};
  assign T17258 = $signed(T17259) / $signed(22'h100000);
  assign T17259 = $signed(30'h28f77ad0) * $signed(16'h1);
  assign T17260 = T17258[6'h2d:6'h2d];
  assign twiddle4_2_317_real = T17263 + T17261;
  assign T17261 = $signed(T17262) / $signed(22'h100000);
  assign T17262 = $signed(31'h3b91af96) * $signed(16'h0);
  assign T17263 = {T17266, T17264};
  assign T17264 = $signed(T17265) / $signed(22'h100000);
  assign T17265 = $signed(30'h2899cbf1) * $signed(16'h1);
  assign T17266 = T17264[6'h2d:6'h2d];
  assign T17267 = T10817[1'h0:1'h0];
  assign T17268 = T17281 ? twiddle4_2_319_real : twiddle4_2_318_real;
  assign twiddle4_2_318_real = T17271 + T17269;
  assign T17269 = $signed(T17270) / $signed(22'h100000);
  assign T17270 = $signed(31'h3b6ca4c4) * $signed(16'h0);
  assign T17271 = {T17274, T17272};
  assign T17272 = $signed(T17273) / $signed(22'h100000);
  assign T17273 = $signed(30'h283c56cf) * $signed(16'h1);
  assign T17274 = T17272[6'h2d:6'h2d];
  assign twiddle4_2_319_real = T17277 + T17275;
  assign T17275 = $signed(T17276) / $signed(22'h100000);
  assign T17276 = $signed(31'h3b470752) * $signed(16'h0);
  assign T17277 = {T17280, T17278};
  assign T17278 = $signed(T17279) / $signed(22'h100000);
  assign T17279 = $signed(30'h27df1c50) * $signed(16'h1);
  assign T17280 = T17278[6'h2d:6'h2d];
  assign T17281 = T10817[1'h0:1'h0];
  assign T17282 = T10817[1'h1:1'h1];
  assign T17283 = T10817[2'h2:2'h2];
  assign T17284 = T10817[2'h3:2'h3];
  assign T17285 = T10817[3'h4:3'h4];
  assign T17286 = T17022[6'h2e:6'h2e];
  assign T17287 = T10817[3'h5:3'h5];
  assign T17288 = {T17715, T17289};
  assign T17289 = T17714 ? T17524 : T17290;
  assign T17290 = T17523 ? T17417 : T17291;
  assign T17291 = T17416 ? T17354 : T17292;
  assign T17292 = T17353 ? T17323 : T17293;
  assign T17293 = T17322 ? T17308 : T17294;
  assign T17294 = T17307 ? twiddle4_2_321_real : twiddle4_2_320_real;
  assign twiddle4_2_320_real = T17297 + T17295;
  assign T17295 = $signed(T17296) / $signed(22'h100000);
  assign T17296 = $signed(31'h3b20d79e) * $signed(16'h0);
  assign T17297 = {T17300, T17298};
  assign T17298 = $signed(T17299) / $signed(22'h100000);
  assign T17299 = $signed(30'h27821d5a) * $signed(16'h1);
  assign T17300 = T17298[6'h2d:6'h2d];
  assign twiddle4_2_321_real = T17303 + T17301;
  assign T17301 = $signed(T17302) / $signed(22'h100000);
  assign T17302 = $signed(31'h3afa1605) * $signed(16'h0);
  assign T17303 = {T17306, T17304};
  assign T17304 = $signed(T17305) / $signed(22'h100000);
  assign T17305 = $signed(30'h27255ad2) * $signed(16'h1);
  assign T17306 = T17304[6'h2d:6'h2d];
  assign T17307 = T10817[1'h0:1'h0];
  assign T17308 = T17321 ? twiddle4_2_323_real : twiddle4_2_322_real;
  assign twiddle4_2_322_real = T17311 + T17309;
  assign T17309 = $signed(T17310) / $signed(22'h100000);
  assign T17310 = $signed(31'h3ad2c2e7) * $signed(16'h0);
  assign T17311 = {T17314, T17312};
  assign T17312 = $signed(T17313) / $signed(22'h100000);
  assign T17313 = $signed(30'h26c8d59d) * $signed(16'h1);
  assign T17314 = T17312[6'h2d:6'h2d];
  assign twiddle4_2_323_real = T17317 + T17315;
  assign T17315 = $signed(T17316) / $signed(22'h100000);
  assign T17316 = $signed(31'h3aaadea5) * $signed(16'h0);
  assign T17317 = {T17320, T17318};
  assign T17318 = $signed(T17319) / $signed(22'h100000);
  assign T17319 = $signed(30'h266c8e9f) * $signed(16'h1);
  assign T17320 = T17318[6'h2d:6'h2d];
  assign T17321 = T10817[1'h0:1'h0];
  assign T17322 = T10817[1'h1:1'h1];
  assign T17323 = T17352 ? T17338 : T17324;
  assign T17324 = T17337 ? twiddle4_2_325_real : twiddle4_2_324_real;
  assign twiddle4_2_324_real = T17327 + T17325;
  assign T17325 = $signed(T17326) / $signed(22'h100000);
  assign T17326 = $signed(31'h3a8269a2) * $signed(16'h0);
  assign T17327 = {T17330, T17328};
  assign T17328 = $signed(T17329) / $signed(22'h100000);
  assign T17329 = $signed(30'h261086bd) * $signed(16'h1);
  assign T17330 = T17328[6'h2d:6'h2d];
  assign twiddle4_2_325_real = T17333 + T17331;
  assign T17331 = $signed(T17332) / $signed(22'h100000);
  assign T17332 = $signed(31'h3a596441) * $signed(16'h0);
  assign T17333 = {T17336, T17334};
  assign T17334 = $signed(T17335) / $signed(22'h100000);
  assign T17335 = $signed(30'h25b4bed9) * $signed(16'h1);
  assign T17336 = T17334[6'h2d:6'h2d];
  assign T17337 = T10817[1'h0:1'h0];
  assign T17338 = T17351 ? twiddle4_2_327_real : twiddle4_2_326_real;
  assign twiddle4_2_326_real = T17341 + T17339;
  assign T17339 = $signed(T17340) / $signed(22'h100000);
  assign T17340 = $signed(31'h3a2fcee8) * $signed(16'h0);
  assign T17341 = {T17344, T17342};
  assign T17342 = $signed(T17343) / $signed(22'h100000);
  assign T17343 = $signed(30'h255937d5) * $signed(16'h1);
  assign T17344 = T17342[6'h2d:6'h2d];
  assign twiddle4_2_327_real = T17347 + T17345;
  assign T17345 = $signed(T17346) / $signed(22'h100000);
  assign T17346 = $signed(31'h3a05a9fd) * $signed(16'h0);
  assign T17347 = {T17350, T17348};
  assign T17348 = $signed(T17349) / $signed(22'h100000);
  assign T17349 = $signed(30'h24fdf294) * $signed(16'h1);
  assign T17350 = T17348[6'h2d:6'h2d];
  assign T17351 = T10817[1'h0:1'h0];
  assign T17352 = T10817[1'h1:1'h1];
  assign T17353 = T10817[2'h2:2'h2];
  assign T17354 = T17415 ? T17385 : T17355;
  assign T17355 = T17384 ? T17370 : T17356;
  assign T17356 = T17369 ? twiddle4_2_329_real : twiddle4_2_328_real;
  assign twiddle4_2_328_real = T17359 + T17357;
  assign T17357 = $signed(T17358) / $signed(22'h100000);
  assign T17358 = $signed(31'h39daf5e8) * $signed(16'h0);
  assign T17359 = {T17362, T17360};
  assign T17360 = $signed(T17361) / $signed(22'h100000);
  assign T17361 = $signed(30'h24a2eff7) * $signed(16'h1);
  assign T17362 = T17360[6'h2d:6'h2d];
  assign twiddle4_2_329_real = T17365 + T17363;
  assign T17363 = $signed(T17364) / $signed(22'h100000);
  assign T17364 = $signed(31'h39afb313) * $signed(16'h0);
  assign T17365 = {T17368, T17366};
  assign T17366 = $signed(T17367) / $signed(22'h100000);
  assign T17367 = $signed(30'h244830dd) * $signed(16'h1);
  assign T17368 = T17366[6'h2d:6'h2d];
  assign T17369 = T10817[1'h0:1'h0];
  assign T17370 = T17383 ? twiddle4_2_331_real : twiddle4_2_330_real;
  assign twiddle4_2_330_real = T17373 + T17371;
  assign T17371 = $signed(T17372) / $signed(22'h100000);
  assign T17372 = $signed(31'h3983e1e7) * $signed(16'h0);
  assign T17373 = {T17376, T17374};
  assign T17374 = $signed(T17375) / $signed(22'h100000);
  assign T17375 = $signed(30'h23edb628) * $signed(16'h1);
  assign T17376 = T17374[6'h2d:6'h2d];
  assign twiddle4_2_331_real = T17379 + T17377;
  assign T17377 = $signed(T17378) / $signed(22'h100000);
  assign T17378 = $signed(31'h395782d3) * $signed(16'h0);
  assign T17379 = {T17382, T17380};
  assign T17380 = $signed(T17381) / $signed(22'h100000);
  assign T17381 = $signed(30'h239380b7) * $signed(16'h1);
  assign T17382 = T17380[6'h2d:6'h2d];
  assign T17383 = T10817[1'h0:1'h0];
  assign T17384 = T10817[1'h1:1'h1];
  assign T17385 = T17414 ? T17400 : T17386;
  assign T17386 = T17399 ? twiddle4_2_333_real : twiddle4_2_332_real;
  assign twiddle4_2_332_real = T17389 + T17387;
  assign T17387 = $signed(T17388) / $signed(22'h100000);
  assign T17388 = $signed(31'h392a9642) * $signed(16'h0);
  assign T17389 = {T17392, T17390};
  assign T17390 = $signed(T17391) / $signed(22'h100000);
  assign T17391 = $signed(30'h23399167) * $signed(16'h1);
  assign T17392 = T17390[6'h2d:6'h2d];
  assign twiddle4_2_333_real = T17395 + T17393;
  assign T17393 = $signed(T17394) / $signed(22'h100000);
  assign T17394 = $signed(31'h38fd1ca4) * $signed(16'h0);
  assign T17395 = {T17398, T17396};
  assign T17396 = $signed(T17397) / $signed(22'h100000);
  assign T17397 = $signed(30'h22dfe918) * $signed(16'h1);
  assign T17398 = T17396[6'h2d:6'h2d];
  assign T17399 = T10817[1'h0:1'h0];
  assign T17400 = T17413 ? twiddle4_2_335_real : twiddle4_2_334_real;
  assign twiddle4_2_334_real = T17403 + T17401;
  assign T17401 = $signed(T17402) / $signed(22'h100000);
  assign T17402 = $signed(31'h38cf1669) * $signed(16'h0);
  assign T17403 = {T17406, T17404};
  assign T17404 = $signed(T17405) / $signed(22'h100000);
  assign T17405 = $signed(30'h228688a5) * $signed(16'h1);
  assign T17406 = T17404[6'h2d:6'h2d];
  assign twiddle4_2_335_real = T17409 + T17407;
  assign T17407 = $signed(T17408) / $signed(22'h100000);
  assign T17408 = $signed(31'h38a08402) * $signed(16'h0);
  assign T17409 = {T17412, T17410};
  assign T17410 = $signed(T17411) / $signed(22'h100000);
  assign T17411 = $signed(30'h222d70ec) * $signed(16'h1);
  assign T17412 = T17410[6'h2d:6'h2d];
  assign T17413 = T10817[1'h0:1'h0];
  assign T17414 = T10817[1'h1:1'h1];
  assign T17415 = T10817[2'h2:2'h2];
  assign T17416 = T10817[2'h3:2'h3];
  assign T17417 = T17522 ? T17476 : T17418;
  assign T17418 = T17475 ? T17449 : T17419;
  assign T17419 = T17448 ? T17434 : T17420;
  assign T17420 = T17433 ? twiddle4_2_337_real : twiddle4_2_336_real;
  assign twiddle4_2_336_real = T17423 + T17421;
  assign T17421 = $signed(T17422) / $signed(22'h100000);
  assign T17422 = $signed(31'h387165e3) * $signed(16'h0);
  assign T17423 = {T17426, T17424};
  assign T17424 = $signed(T17425) / $signed(22'h100000);
  assign T17425 = $signed(30'h21d4a2c8) * $signed(16'h1);
  assign T17426 = T17424[6'h2d:6'h2d];
  assign twiddle4_2_337_real = T17429 + T17427;
  assign T17427 = $signed(T17428) / $signed(22'h100000);
  assign T17428 = $signed(31'h3841bc7f) * $signed(16'h0);
  assign T17429 = {T17432, T17430};
  assign T17430 = $signed(T17431) / $signed(22'h100000);
  assign T17431 = $signed(30'h217c1f16) * $signed(16'h1);
  assign T17432 = T17430[6'h2d:6'h2d];
  assign T17433 = T10817[1'h0:1'h0];
  assign T17434 = T17447 ? twiddle4_2_339_real : twiddle4_2_338_real;
  assign twiddle4_2_338_real = T17437 + T17435;
  assign T17435 = $signed(T17436) / $signed(22'h100000);
  assign T17436 = $signed(31'h3811884c) * $signed(16'h0);
  assign T17437 = {T17440, T17438};
  assign T17438 = $signed(T17439) / $signed(22'h100000);
  assign T17439 = $signed(30'h2123e6ae) * $signed(16'h1);
  assign T17440 = T17438[6'h2d:6'h2d];
  assign twiddle4_2_339_real = T17443 + T17441;
  assign T17441 = $signed(T17442) / $signed(22'h100000);
  assign T17442 = $signed(31'h37e0c9c2) * $signed(16'h0);
  assign T17443 = {T17446, T17444};
  assign T17444 = $signed(T17445) / $signed(22'h100000);
  assign T17445 = $signed(30'h20cbfa6a) * $signed(16'h1);
  assign T17446 = T17444[6'h2d:6'h2d];
  assign T17447 = T10817[1'h0:1'h0];
  assign T17448 = T10817[1'h1:1'h1];
  assign T17449 = T17474 ? T17464 : T17450;
  assign T17450 = T17463 ? twiddle4_2_341_real : twiddle4_2_340_real;
  assign twiddle4_2_340_real = T17453 + T17451;
  assign T17451 = $signed(T17452) / $signed(22'h100000);
  assign T17452 = $signed(31'h37af8158) * $signed(16'h0);
  assign T17453 = {T17456, T17454};
  assign T17454 = $signed(T17455) / $signed(22'h100000);
  assign T17455 = $signed(30'h20745b25) * $signed(16'h1);
  assign T17456 = T17454[6'h2d:6'h2d];
  assign twiddle4_2_341_real = T17459 + T17457;
  assign T17457 = $signed(T17458) / $signed(22'h100000);
  assign T17458 = $signed(31'h377daf89) * $signed(16'h0);
  assign T17459 = {T17462, T17460};
  assign T17460 = $signed(T17461) / $signed(22'h100000);
  assign T17461 = $signed(30'h201d09b5) * $signed(16'h1);
  assign T17462 = T17460[6'h2d:6'h2d];
  assign T17463 = T10817[1'h0:1'h0];
  assign T17464 = T17473 ? twiddle4_2_343_real : twiddle4_2_342_real;
  assign twiddle4_2_342_real = T17467 + T17465;
  assign T17465 = $signed(T17466) / $signed(22'h100000);
  assign T17466 = $signed(31'h374b54ce) * $signed(16'h0);
  assign T17467 = $signed(T17468) / $signed(22'h100000);
  assign T17468 = $signed(31'h5fc606f2) * $signed(16'h1);
  assign twiddle4_2_343_real = T17471 + T17469;
  assign T17469 = $signed(T17470) / $signed(22'h100000);
  assign T17470 = $signed(31'h371871a4) * $signed(16'h0);
  assign T17471 = $signed(T17472) / $signed(22'h100000);
  assign T17472 = $signed(31'h5f6f53b3) * $signed(16'h1);
  assign T17473 = T10817[1'h0:1'h0];
  assign T17474 = T10817[1'h1:1'h1];
  assign T17475 = T10817[2'h2:2'h2];
  assign T17476 = T17521 ? T17499 : T17477;
  assign T17477 = T17498 ? T17488 : T17478;
  assign T17478 = T17487 ? twiddle4_2_345_real : twiddle4_2_344_real;
  assign twiddle4_2_344_real = T17481 + T17479;
  assign T17479 = $signed(T17480) / $signed(22'h100000);
  assign T17480 = $signed(31'h36e5068a) * $signed(16'h0);
  assign T17481 = $signed(T17482) / $signed(22'h100000);
  assign T17482 = $signed(31'h5f18f0ce) * $signed(16'h1);
  assign twiddle4_2_345_real = T17485 + T17483;
  assign T17483 = $signed(T17484) / $signed(22'h100000);
  assign T17484 = $signed(31'h36b113fd) * $signed(16'h0);
  assign T17485 = $signed(T17486) / $signed(22'h100000);
  assign T17486 = $signed(31'h5ec2df18) * $signed(16'h1);
  assign T17487 = T10817[1'h0:1'h0];
  assign T17488 = T17497 ? twiddle4_2_347_real : twiddle4_2_346_real;
  assign twiddle4_2_346_real = T17491 + T17489;
  assign T17489 = $signed(T17490) / $signed(22'h100000);
  assign T17490 = $signed(31'h367c9a7d) * $signed(16'h0);
  assign T17491 = $signed(T17492) / $signed(22'h100000);
  assign T17492 = $signed(31'h5e6d1f66) * $signed(16'h1);
  assign twiddle4_2_347_real = T17495 + T17493;
  assign T17493 = $signed(T17494) / $signed(22'h100000);
  assign T17494 = $signed(31'h36479a8e) * $signed(16'h0);
  assign T17495 = $signed(T17496) / $signed(22'h100000);
  assign T17496 = $signed(31'h5e17b28a) * $signed(16'h1);
  assign T17497 = T10817[1'h0:1'h0];
  assign T17498 = T10817[1'h1:1'h1];
  assign T17499 = T17520 ? T17510 : T17500;
  assign T17500 = T17509 ? twiddle4_2_349_real : twiddle4_2_348_real;
  assign twiddle4_2_348_real = T17503 + T17501;
  assign T17501 = $signed(T17502) / $signed(22'h100000);
  assign T17502 = $signed(31'h361214b0) * $signed(16'h0);
  assign T17503 = $signed(T17504) / $signed(22'h100000);
  assign T17504 = $signed(31'h5dc29958) * $signed(16'h1);
  assign twiddle4_2_349_real = T17507 + T17505;
  assign T17505 = $signed(T17506) / $signed(22'h100000);
  assign T17506 = $signed(31'h35dc0968) * $signed(16'h0);
  assign T17507 = $signed(T17508) / $signed(22'h100000);
  assign T17508 = $signed(31'h5d6dd4a2) * $signed(16'h1);
  assign T17509 = T10817[1'h0:1'h0];
  assign T17510 = T17519 ? twiddle4_2_351_real : twiddle4_2_350_real;
  assign twiddle4_2_350_real = T17513 + T17511;
  assign T17511 = $signed(T17512) / $signed(22'h100000);
  assign T17512 = $signed(31'h35a5793c) * $signed(16'h0);
  assign T17513 = $signed(T17514) / $signed(22'h100000);
  assign T17514 = $signed(31'h5d196539) * $signed(16'h1);
  assign twiddle4_2_351_real = T17517 + T17515;
  assign T17515 = $signed(T17516) / $signed(22'h100000);
  assign T17516 = $signed(31'h356e64b2) * $signed(16'h0);
  assign T17517 = $signed(T17518) / $signed(22'h100000);
  assign T17518 = $signed(31'h5cc54bed) * $signed(16'h1);
  assign T17519 = T10817[1'h0:1'h0];
  assign T17520 = T10817[1'h1:1'h1];
  assign T17521 = T10817[2'h2:2'h2];
  assign T17522 = T10817[2'h3:2'h3];
  assign T17523 = T10817[3'h4:3'h4];
  assign T17524 = T17713 ? T17619 : T17525;
  assign T17525 = T17618 ? T17572 : T17526;
  assign T17526 = T17571 ? T17549 : T17527;
  assign T17527 = T17548 ? T17538 : T17528;
  assign T17528 = T17537 ? twiddle4_2_353_real : twiddle4_2_352_real;
  assign twiddle4_2_352_real = T17531 + T17529;
  assign T17529 = $signed(T17530) / $signed(22'h100000);
  assign T17530 = $signed(31'h3536cc52) * $signed(16'h0);
  assign T17531 = $signed(T17532) / $signed(22'h100000);
  assign T17532 = $signed(31'h5c71898d) * $signed(16'h1);
  assign twiddle4_2_353_real = T17535 + T17533;
  assign T17533 = $signed(T17534) / $signed(22'h100000);
  assign T17534 = $signed(31'h34feb0a5) * $signed(16'h0);
  assign T17535 = $signed(T17536) / $signed(22'h100000);
  assign T17536 = $signed(31'h5c1e1ee9) * $signed(16'h1);
  assign T17537 = T10817[1'h0:1'h0];
  assign T17538 = T17547 ? twiddle4_2_355_real : twiddle4_2_354_real;
  assign twiddle4_2_354_real = T17541 + T17539;
  assign T17539 = $signed(T17540) / $signed(22'h100000);
  assign T17540 = $signed(31'h34c61236) * $signed(16'h0);
  assign T17541 = $signed(T17542) / $signed(22'h100000);
  assign T17542 = $signed(31'h5bcb0cce) * $signed(16'h1);
  assign twiddle4_2_355_real = T17545 + T17543;
  assign T17543 = $signed(T17544) / $signed(22'h100000);
  assign T17544 = $signed(31'h348cf190) * $signed(16'h0);
  assign T17545 = $signed(T17546) / $signed(22'h100000);
  assign T17546 = $signed(31'h5b785409) * $signed(16'h1);
  assign T17547 = T10817[1'h0:1'h0];
  assign T17548 = T10817[1'h1:1'h1];
  assign T17549 = T17570 ? T17560 : T17550;
  assign T17550 = T17559 ? twiddle4_2_357_real : twiddle4_2_356_real;
  assign twiddle4_2_356_real = T17553 + T17551;
  assign T17551 = $signed(T17552) / $signed(22'h100000);
  assign T17552 = $signed(31'h34534f40) * $signed(16'h0);
  assign T17553 = $signed(T17554) / $signed(22'h100000);
  assign T17554 = $signed(31'h5b25f567) * $signed(16'h1);
  assign twiddle4_2_357_real = T17557 + T17555;
  assign T17555 = $signed(T17556) / $signed(22'h100000);
  assign T17556 = $signed(31'h34192bd5) * $signed(16'h0);
  assign T17557 = $signed(T17558) / $signed(22'h100000);
  assign T17558 = $signed(31'h5ad3f1b2) * $signed(16'h1);
  assign T17559 = T10817[1'h0:1'h0];
  assign T17560 = T17569 ? twiddle4_2_359_real : twiddle4_2_358_real;
  assign twiddle4_2_358_real = T17563 + T17561;
  assign T17561 = $signed(T17562) / $signed(22'h100000);
  assign T17562 = $signed(31'h33de87de) * $signed(16'h0);
  assign T17563 = $signed(T17564) / $signed(22'h100000);
  assign T17564 = $signed(31'h5a8249b5) * $signed(16'h1);
  assign twiddle4_2_359_real = T17567 + T17565;
  assign T17565 = $signed(T17566) / $signed(22'h100000);
  assign T17566 = $signed(31'h33a363eb) * $signed(16'h0);
  assign T17567 = $signed(T17568) / $signed(22'h100000);
  assign T17568 = $signed(31'h5a30fe39) * $signed(16'h1);
  assign T17569 = T10817[1'h0:1'h0];
  assign T17570 = T10817[1'h1:1'h1];
  assign T17571 = T10817[2'h2:2'h2];
  assign T17572 = T17617 ? T17595 : T17573;
  assign T17573 = T17594 ? T17584 : T17574;
  assign T17574 = T17583 ? twiddle4_2_361_real : twiddle4_2_360_real;
  assign twiddle4_2_360_real = T17577 + T17575;
  assign T17575 = $signed(T17576) / $signed(22'h100000);
  assign T17576 = $signed(31'h3367c08f) * $signed(16'h0);
  assign T17577 = $signed(T17578) / $signed(22'h100000);
  assign T17578 = $signed(31'h59e01007) * $signed(16'h1);
  assign twiddle4_2_361_real = T17581 + T17579;
  assign T17579 = $signed(T17580) / $signed(22'h100000);
  assign T17580 = $signed(31'h332b9e5d) * $signed(16'h0);
  assign T17581 = $signed(T17582) / $signed(22'h100000);
  assign T17582 = $signed(31'h598f7fe6) * $signed(16'h1);
  assign T17583 = T10817[1'h0:1'h0];
  assign T17584 = T17593 ? twiddle4_2_363_real : twiddle4_2_362_real;
  assign twiddle4_2_362_real = T17587 + T17585;
  assign T17585 = $signed(T17586) / $signed(22'h100000);
  assign T17586 = $signed(31'h32eefde9) * $signed(16'h0);
  assign T17587 = $signed(T17588) / $signed(22'h100000);
  assign T17588 = $signed(31'h593f4e9e) * $signed(16'h1);
  assign twiddle4_2_363_real = T17591 + T17589;
  assign T17589 = $signed(T17590) / $signed(22'h100000);
  assign T17590 = $signed(31'h32b1dfc9) * $signed(16'h0);
  assign T17591 = $signed(T17592) / $signed(22'h100000);
  assign T17592 = $signed(31'h58ef7cf5) * $signed(16'h1);
  assign T17593 = T10817[1'h0:1'h0];
  assign T17594 = T10817[1'h1:1'h1];
  assign T17595 = T17616 ? T17606 : T17596;
  assign T17596 = T17605 ? twiddle4_2_365_real : twiddle4_2_364_real;
  assign twiddle4_2_364_real = T17599 + T17597;
  assign T17597 = $signed(T17598) / $signed(22'h100000);
  assign T17598 = $signed(31'h32744493) * $signed(16'h0);
  assign T17599 = $signed(T17600) / $signed(22'h100000);
  assign T17600 = $signed(31'h58a00bae) * $signed(16'h1);
  assign twiddle4_2_365_real = T17603 + T17601;
  assign T17601 = $signed(T17602) / $signed(22'h100000);
  assign T17602 = $signed(31'h32362cdf) * $signed(16'h0);
  assign T17603 = $signed(T17604) / $signed(22'h100000);
  assign T17604 = $signed(31'h5850fb8f) * $signed(16'h1);
  assign T17605 = T10817[1'h0:1'h0];
  assign T17606 = T17615 ? twiddle4_2_367_real : twiddle4_2_366_real;
  assign twiddle4_2_366_real = T17609 + T17607;
  assign T17607 = $signed(T17608) / $signed(22'h100000);
  assign T17608 = $signed(31'h31f79947) * $signed(16'h0);
  assign T17609 = $signed(T17610) / $signed(22'h100000);
  assign T17610 = $signed(31'h58024d5a) * $signed(16'h1);
  assign twiddle4_2_367_real = T17613 + T17611;
  assign T17611 = $signed(T17612) / $signed(22'h100000);
  assign T17612 = $signed(31'h31b88a66) * $signed(16'h0);
  assign T17613 = $signed(T17614) / $signed(22'h100000);
  assign T17614 = $signed(31'h57b401d1) * $signed(16'h1);
  assign T17615 = T10817[1'h0:1'h0];
  assign T17616 = T10817[1'h1:1'h1];
  assign T17617 = T10817[2'h2:2'h2];
  assign T17618 = T10817[2'h3:2'h3];
  assign T17619 = T17712 ? T17666 : T17620;
  assign T17620 = T17665 ? T17643 : T17621;
  assign T17621 = T17642 ? T17632 : T17622;
  assign T17622 = T17631 ? twiddle4_2_369_real : twiddle4_2_368_real;
  assign twiddle4_2_368_real = T17625 + T17623;
  assign T17623 = $signed(T17624) / $signed(22'h100000);
  assign T17624 = $signed(31'h317900d6) * $signed(16'h0);
  assign T17625 = $signed(T17626) / $signed(22'h100000);
  assign T17626 = $signed(31'h576619b6) * $signed(16'h1);
  assign twiddle4_2_369_real = T17629 + T17627;
  assign T17627 = $signed(T17628) / $signed(22'h100000);
  assign T17628 = $signed(31'h3138fd34) * $signed(16'h0);
  assign T17629 = $signed(T17630) / $signed(22'h100000);
  assign T17630 = $signed(31'h571895c9) * $signed(16'h1);
  assign T17631 = T10817[1'h0:1'h0];
  assign T17632 = T17641 ? twiddle4_2_371_real : twiddle4_2_370_real;
  assign twiddle4_2_370_real = T17635 + T17633;
  assign T17633 = $signed(T17634) / $signed(22'h100000);
  assign T17634 = $signed(31'h30f8801f) * $signed(16'h0);
  assign T17635 = $signed(T17636) / $signed(22'h100000);
  assign T17636 = $signed(31'h56cb76c9) * $signed(16'h1);
  assign twiddle4_2_371_real = T17639 + T17637;
  assign T17637 = $signed(T17638) / $signed(22'h100000);
  assign T17638 = $signed(31'h30b78a35) * $signed(16'h0);
  assign T17639 = $signed(T17640) / $signed(22'h100000);
  assign T17640 = $signed(31'h567ebd75) * $signed(16'h1);
  assign T17641 = T10817[1'h0:1'h0];
  assign T17642 = T10817[1'h1:1'h1];
  assign T17643 = T17664 ? T17654 : T17644;
  assign T17644 = T17653 ? twiddle4_2_373_real : twiddle4_2_372_real;
  assign twiddle4_2_372_real = T17647 + T17645;
  assign T17645 = $signed(T17646) / $signed(22'h100000);
  assign T17646 = $signed(31'h30761c17) * $signed(16'h0);
  assign T17647 = $signed(T17648) / $signed(22'h100000);
  assign T17648 = $signed(31'h56326a89) * $signed(16'h1);
  assign twiddle4_2_373_real = T17651 + T17649;
  assign T17649 = $signed(T17650) / $signed(22'h100000);
  assign T17650 = $signed(31'h30343667) * $signed(16'h0);
  assign T17651 = $signed(T17652) / $signed(22'h100000);
  assign T17652 = $signed(31'h55e67ec2) * $signed(16'h1);
  assign T17653 = T10817[1'h0:1'h0];
  assign T17654 = T17663 ? twiddle4_2_375_real : twiddle4_2_374_real;
  assign twiddle4_2_374_real = T17657 + T17655;
  assign T17655 = $signed(T17656) / $signed(22'h100000);
  assign T17656 = $signed(31'h2ff1d9c6) * $signed(16'h0);
  assign T17657 = $signed(T17658) / $signed(22'h100000);
  assign T17658 = $signed(31'h559afadb) * $signed(16'h1);
  assign twiddle4_2_375_real = T17661 + T17659;
  assign T17659 = $signed(T17660) / $signed(22'h100000);
  assign T17660 = $signed(31'h2faf06d9) * $signed(16'h0);
  assign T17661 = $signed(T17662) / $signed(22'h100000);
  assign T17662 = $signed(31'h554fdf8f) * $signed(16'h1);
  assign T17663 = T10817[1'h0:1'h0];
  assign T17664 = T10817[1'h1:1'h1];
  assign T17665 = T10817[2'h2:2'h2];
  assign T17666 = T17711 ? T17689 : T17667;
  assign T17667 = T17688 ? T17678 : T17668;
  assign T17668 = T17677 ? twiddle4_2_377_real : twiddle4_2_376_real;
  assign twiddle4_2_376_real = T17671 + T17669;
  assign T17669 = $signed(T17670) / $signed(22'h100000);
  assign T17670 = $signed(31'h2f6bbe44) * $signed(16'h0);
  assign T17671 = $signed(T17672) / $signed(22'h100000);
  assign T17672 = $signed(31'h55052d97) * $signed(16'h1);
  assign twiddle4_2_377_real = T17675 + T17673;
  assign T17673 = $signed(T17674) / $signed(22'h100000);
  assign T17674 = $signed(31'h2f2800ae) * $signed(16'h0);
  assign T17675 = $signed(T17676) / $signed(22'h100000);
  assign T17676 = $signed(31'h54bae5ac) * $signed(16'h1);
  assign T17677 = T10817[1'h0:1'h0];
  assign T17678 = T17687 ? twiddle4_2_379_real : twiddle4_2_378_real;
  assign twiddle4_2_378_real = T17681 + T17679;
  assign T17679 = $signed(T17680) / $signed(22'h100000);
  assign T17680 = $signed(31'h2ee3cebe) * $signed(16'h0);
  assign T17681 = $signed(T17682) / $signed(22'h100000);
  assign T17682 = $signed(31'h54710884) * $signed(16'h1);
  assign twiddle4_2_379_real = T17685 + T17683;
  assign T17683 = $signed(T17684) / $signed(22'h100000);
  assign T17684 = $signed(31'h2e9f291b) * $signed(16'h0);
  assign T17685 = $signed(T17686) / $signed(22'h100000);
  assign T17686 = $signed(31'h542796d5) * $signed(16'h1);
  assign T17687 = T10817[1'h0:1'h0];
  assign T17688 = T10817[1'h1:1'h1];
  assign T17689 = T17710 ? T17700 : T17690;
  assign T17690 = T17699 ? twiddle4_2_381_real : twiddle4_2_380_real;
  assign twiddle4_2_380_real = T17693 + T17691;
  assign T17691 = $signed(T17692) / $signed(22'h100000);
  assign T17692 = $signed(31'h2e5a106f) * $signed(16'h0);
  assign T17693 = $signed(T17694) / $signed(22'h100000);
  assign T17694 = $signed(31'h53de9156) * $signed(16'h1);
  assign twiddle4_2_381_real = T17697 + T17695;
  assign T17695 = $signed(T17696) / $signed(22'h100000);
  assign T17696 = $signed(31'h2e148566) * $signed(16'h0);
  assign T17697 = $signed(T17698) / $signed(22'h100000);
  assign T17698 = $signed(31'h5395f8ba) * $signed(16'h1);
  assign T17699 = T10817[1'h0:1'h0];
  assign T17700 = T17709 ? twiddle4_2_383_real : twiddle4_2_382_real;
  assign twiddle4_2_382_real = T17703 + T17701;
  assign T17701 = $signed(T17702) / $signed(22'h100000);
  assign T17702 = $signed(31'h2dce88a9) * $signed(16'h0);
  assign T17703 = $signed(T17704) / $signed(22'h100000);
  assign T17704 = $signed(31'h534dcdb5) * $signed(16'h1);
  assign twiddle4_2_383_real = T17707 + T17705;
  assign T17705 = $signed(T17706) / $signed(22'h100000);
  assign T17706 = $signed(31'h2d881ae7) * $signed(16'h0);
  assign T17707 = $signed(T17708) / $signed(22'h100000);
  assign T17708 = $signed(31'h530610f7) * $signed(16'h1);
  assign T17709 = T10817[1'h0:1'h0];
  assign T17710 = T10817[1'h1:1'h1];
  assign T17711 = T10817[2'h2:2'h2];
  assign T17712 = T10817[2'h3:2'h3];
  assign T17713 = T10817[3'h4:3'h4];
  assign T17714 = T10817[3'h5:3'h5];
  assign T17715 = T17289[6'h2e:6'h2e];
  assign T17716 = T10817[3'h6:3'h6];
  assign T17717 = {T18695, T17718};
  assign T17718 = T18694 ? T18143 : T17719;
  assign T17719 = T18142 ? T17910 : T17720;
  assign T17720 = T17909 ? T17815 : T17721;
  assign T17721 = T17814 ? T17768 : T17722;
  assign T17722 = T17767 ? T17745 : T17723;
  assign T17723 = T17744 ? T17734 : T17724;
  assign T17724 = T17733 ? twiddle4_2_385_real : twiddle4_2_384_real;
  assign twiddle4_2_384_real = T17727 + T17725;
  assign T17725 = $signed(T17726) / $signed(22'h100000);
  assign T17726 = $signed(31'h2d413ccc) * $signed(16'h0);
  assign T17727 = $signed(T17728) / $signed(22'h100000);
  assign T17728 = $signed(31'h52bec334) * $signed(16'h1);
  assign twiddle4_2_385_real = T17731 + T17729;
  assign T17729 = $signed(T17730) / $signed(22'h100000);
  assign T17730 = $signed(31'h2cf9ef09) * $signed(16'h0);
  assign T17731 = $signed(T17732) / $signed(22'h100000);
  assign T17732 = $signed(31'h5277e519) * $signed(16'h1);
  assign T17733 = T10817[1'h0:1'h0];
  assign T17734 = T17743 ? twiddle4_2_387_real : twiddle4_2_386_real;
  assign twiddle4_2_386_real = T17737 + T17735;
  assign T17735 = $signed(T17736) / $signed(22'h100000);
  assign T17736 = $signed(31'h2cb2324b) * $signed(16'h0);
  assign T17737 = $signed(T17738) / $signed(22'h100000);
  assign T17738 = $signed(31'h52317757) * $signed(16'h1);
  assign twiddle4_2_387_real = T17741 + T17739;
  assign T17739 = $signed(T17740) / $signed(22'h100000);
  assign T17740 = $signed(31'h2c6a0746) * $signed(16'h0);
  assign T17741 = $signed(T17742) / $signed(22'h100000);
  assign T17742 = $signed(31'h51eb7a9a) * $signed(16'h1);
  assign T17743 = T10817[1'h0:1'h0];
  assign T17744 = T10817[1'h1:1'h1];
  assign T17745 = T17766 ? T17756 : T17746;
  assign T17746 = T17755 ? twiddle4_2_389_real : twiddle4_2_388_real;
  assign twiddle4_2_388_real = T17749 + T17747;
  assign T17747 = $signed(T17748) / $signed(22'h100000);
  assign T17748 = $signed(31'h2c216eaa) * $signed(16'h0);
  assign T17749 = $signed(T17750) / $signed(22'h100000);
  assign T17750 = $signed(31'h51a5ef91) * $signed(16'h1);
  assign twiddle4_2_389_real = T17753 + T17751;
  assign T17751 = $signed(T17752) / $signed(22'h100000);
  assign T17752 = $signed(31'h2bd8692b) * $signed(16'h0);
  assign T17753 = $signed(T17754) / $signed(22'h100000);
  assign T17754 = $signed(31'h5160d6e5) * $signed(16'h1);
  assign T17755 = T10817[1'h0:1'h0];
  assign T17756 = T17765 ? twiddle4_2_391_real : twiddle4_2_390_real;
  assign twiddle4_2_390_real = T17759 + T17757;
  assign T17757 = $signed(T17758) / $signed(22'h100000);
  assign T17758 = $signed(31'h2b8ef77c) * $signed(16'h0);
  assign T17759 = $signed(T17760) / $signed(22'h100000);
  assign T17760 = $signed(31'h511c3142) * $signed(16'h1);
  assign twiddle4_2_391_real = T17763 + T17761;
  assign T17761 = $signed(T17762) / $signed(22'h100000);
  assign T17762 = $signed(31'h2b451a54) * $signed(16'h0);
  assign T17763 = $signed(T17764) / $signed(22'h100000);
  assign T17764 = $signed(31'h50d7ff52) * $signed(16'h1);
  assign T17765 = T10817[1'h0:1'h0];
  assign T17766 = T10817[1'h1:1'h1];
  assign T17767 = T10817[2'h2:2'h2];
  assign T17768 = T17813 ? T17791 : T17769;
  assign T17769 = T17790 ? T17780 : T17770;
  assign T17770 = T17779 ? twiddle4_2_393_real : twiddle4_2_392_real;
  assign twiddle4_2_392_real = T17773 + T17771;
  assign T17771 = $signed(T17772) / $signed(22'h100000);
  assign T17772 = $signed(31'h2afad269) * $signed(16'h0);
  assign T17773 = $signed(T17774) / $signed(22'h100000);
  assign T17774 = $signed(31'h509441bc) * $signed(16'h1);
  assign twiddle4_2_393_real = T17777 + T17775;
  assign T17775 = $signed(T17776) / $signed(22'h100000);
  assign T17776 = $signed(31'h2ab02071) * $signed(16'h0);
  assign T17777 = $signed(T17778) / $signed(22'h100000);
  assign T17778 = $signed(31'h5050f927) * $signed(16'h1);
  assign T17779 = T10817[1'h0:1'h0];
  assign T17780 = T17789 ? twiddle4_2_395_real : twiddle4_2_394_real;
  assign twiddle4_2_394_real = T17783 + T17781;
  assign T17781 = $signed(T17782) / $signed(22'h100000);
  assign T17782 = $signed(31'h2a650525) * $signed(16'h0);
  assign T17783 = $signed(T17784) / $signed(22'h100000);
  assign T17784 = $signed(31'h500e263a) * $signed(16'h1);
  assign twiddle4_2_395_real = T17787 + T17785;
  assign T17785 = $signed(T17786) / $signed(22'h100000);
  assign T17786 = $signed(31'h2a19813e) * $signed(16'h0);
  assign T17787 = $signed(T17788) / $signed(22'h100000);
  assign T17788 = $signed(31'h4fcbc999) * $signed(16'h1);
  assign T17789 = T10817[1'h0:1'h0];
  assign T17790 = T10817[1'h1:1'h1];
  assign T17791 = T17812 ? T17802 : T17792;
  assign T17792 = T17801 ? twiddle4_2_397_real : twiddle4_2_396_real;
  assign twiddle4_2_396_real = T17795 + T17793;
  assign T17793 = $signed(T17794) / $signed(22'h100000);
  assign T17794 = $signed(31'h29cd9577) * $signed(16'h0);
  assign T17795 = $signed(T17796) / $signed(22'h100000);
  assign T17796 = $signed(31'h4f89e3e9) * $signed(16'h1);
  assign twiddle4_2_397_real = T17799 + T17797;
  assign T17797 = $signed(T17798) / $signed(22'h100000);
  assign T17798 = $signed(31'h2981428b) * $signed(16'h0);
  assign T17799 = $signed(T17800) / $signed(22'h100000);
  assign T17800 = $signed(31'h4f4875cb) * $signed(16'h1);
  assign T17801 = T10817[1'h0:1'h0];
  assign T17802 = T17811 ? twiddle4_2_399_real : twiddle4_2_398_real;
  assign twiddle4_2_398_real = T17805 + T17803;
  assign T17803 = $signed(T17804) / $signed(22'h100000);
  assign T17804 = $signed(31'h29348937) * $signed(16'h0);
  assign T17805 = $signed(T17806) / $signed(22'h100000);
  assign T17806 = $signed(31'h4f077fe1) * $signed(16'h1);
  assign twiddle4_2_399_real = T17809 + T17807;
  assign T17807 = $signed(T17808) / $signed(22'h100000);
  assign T17808 = $signed(31'h28e76a37) * $signed(16'h0);
  assign T17809 = $signed(T17810) / $signed(22'h100000);
  assign T17810 = $signed(31'h4ec702cc) * $signed(16'h1);
  assign T17811 = T10817[1'h0:1'h0];
  assign T17812 = T10817[1'h1:1'h1];
  assign T17813 = T10817[2'h2:2'h2];
  assign T17814 = T10817[2'h3:2'h3];
  assign T17815 = T17908 ? T17862 : T17816;
  assign T17816 = T17861 ? T17839 : T17817;
  assign T17817 = T17838 ? T17828 : T17818;
  assign T17818 = T17827 ? twiddle4_2_401_real : twiddle4_2_400_real;
  assign twiddle4_2_400_real = T17821 + T17819;
  assign T17819 = $signed(T17820) / $signed(22'h100000);
  assign T17820 = $signed(31'h2899e64a) * $signed(16'h0);
  assign T17821 = $signed(T17822) / $signed(22'h100000);
  assign T17822 = $signed(31'h4e86ff2a) * $signed(16'h1);
  assign twiddle4_2_401_real = T17825 + T17823;
  assign T17823 = $signed(T17824) / $signed(22'h100000);
  assign T17824 = $signed(31'h284bfe2f) * $signed(16'h0);
  assign T17825 = $signed(T17826) / $signed(22'h100000);
  assign T17826 = $signed(31'h4e47759a) * $signed(16'h1);
  assign T17827 = T10817[1'h0:1'h0];
  assign T17828 = T17837 ? twiddle4_2_403_real : twiddle4_2_402_real;
  assign twiddle4_2_402_real = T17831 + T17829;
  assign T17829 = $signed(T17830) / $signed(22'h100000);
  assign T17830 = $signed(31'h27fdb2a6) * $signed(16'h0);
  assign T17831 = $signed(T17832) / $signed(22'h100000);
  assign T17832 = $signed(31'h4e0866b9) * $signed(16'h1);
  assign twiddle4_2_403_real = T17835 + T17833;
  assign T17833 = $signed(T17834) / $signed(22'h100000);
  assign T17834 = $signed(31'h27af0471) * $signed(16'h0);
  assign T17835 = $signed(T17836) / $signed(22'h100000);
  assign T17836 = $signed(31'h4dc9d321) * $signed(16'h1);
  assign T17837 = T10817[1'h0:1'h0];
  assign T17838 = T10817[1'h1:1'h1];
  assign T17839 = T17860 ? T17850 : T17840;
  assign T17840 = T17849 ? twiddle4_2_405_real : twiddle4_2_404_real;
  assign twiddle4_2_404_real = T17843 + T17841;
  assign T17841 = $signed(T17842) / $signed(22'h100000);
  assign T17842 = $signed(31'h275ff452) * $signed(16'h0);
  assign T17843 = $signed(T17844) / $signed(22'h100000);
  assign T17844 = $signed(31'h4d8bbb6d) * $signed(16'h1);
  assign twiddle4_2_405_real = T17847 + T17845;
  assign T17845 = $signed(T17846) / $signed(22'h100000);
  assign T17846 = $signed(31'h2710830b) * $signed(16'h0);
  assign T17847 = $signed(T17848) / $signed(22'h100000);
  assign T17848 = $signed(31'h4d4e2037) * $signed(16'h1);
  assign T17849 = T10817[1'h0:1'h0];
  assign T17850 = T17859 ? twiddle4_2_407_real : twiddle4_2_406_real;
  assign twiddle4_2_406_real = T17853 + T17851;
  assign T17851 = $signed(T17852) / $signed(22'h100000);
  assign T17852 = $signed(31'h26c0b162) * $signed(16'h0);
  assign T17853 = $signed(T17854) / $signed(22'h100000);
  assign T17854 = $signed(31'h4d110217) * $signed(16'h1);
  assign twiddle4_2_407_real = T17857 + T17855;
  assign T17855 = $signed(T17856) / $signed(22'h100000);
  assign T17856 = $signed(31'h2670801a) * $signed(16'h0);
  assign T17857 = $signed(T17858) / $signed(22'h100000);
  assign T17858 = $signed(31'h4cd461a3) * $signed(16'h1);
  assign T17859 = T10817[1'h0:1'h0];
  assign T17860 = T10817[1'h1:1'h1];
  assign T17861 = T10817[2'h2:2'h2];
  assign T17862 = T17907 ? T17885 : T17863;
  assign T17863 = T17884 ? T17874 : T17864;
  assign T17864 = T17873 ? twiddle4_2_409_real : twiddle4_2_408_real;
  assign twiddle4_2_408_real = T17867 + T17865;
  assign T17865 = $signed(T17866) / $signed(22'h100000);
  assign T17866 = $signed(31'h261feff9) * $signed(16'h0);
  assign T17867 = $signed(T17868) / $signed(22'h100000);
  assign T17868 = $signed(31'h4c983f71) * $signed(16'h1);
  assign twiddle4_2_409_real = T17871 + T17869;
  assign T17869 = $signed(T17870) / $signed(22'h100000);
  assign T17870 = $signed(31'h25cf01c7) * $signed(16'h0);
  assign T17871 = $signed(T17872) / $signed(22'h100000);
  assign T17872 = $signed(31'h4c5c9c15) * $signed(16'h1);
  assign T17873 = T10817[1'h0:1'h0];
  assign T17874 = T17883 ? twiddle4_2_411_real : twiddle4_2_410_real;
  assign twiddle4_2_410_real = T17877 + T17875;
  assign T17875 = $signed(T17876) / $signed(22'h100000);
  assign T17876 = $signed(31'h257db64b) * $signed(16'h0);
  assign T17877 = $signed(T17878) / $signed(22'h100000);
  assign T17878 = $signed(31'h4c217822) * $signed(16'h1);
  assign twiddle4_2_411_real = T17881 + T17879;
  assign T17879 = $signed(T17880) / $signed(22'h100000);
  assign T17880 = $signed(31'h252c0e4e) * $signed(16'h0);
  assign T17881 = $signed(T17882) / $signed(22'h100000);
  assign T17882 = $signed(31'h4be6d42b) * $signed(16'h1);
  assign T17883 = T10817[1'h0:1'h0];
  assign T17884 = T10817[1'h1:1'h1];
  assign T17885 = T17906 ? T17896 : T17886;
  assign T17886 = T17895 ? twiddle4_2_413_real : twiddle4_2_412_real;
  assign twiddle4_2_412_real = T17889 + T17887;
  assign T17887 = $signed(T17888) / $signed(22'h100000);
  assign T17888 = $signed(31'h24da0a99) * $signed(16'h0);
  assign T17889 = $signed(T17890) / $signed(22'h100000);
  assign T17890 = $signed(31'h4bacb0c0) * $signed(16'h1);
  assign twiddle4_2_413_real = T17893 + T17891;
  assign T17891 = $signed(T17892) / $signed(22'h100000);
  assign T17892 = $signed(31'h2487abf7) * $signed(16'h0);
  assign T17893 = $signed(T17894) / $signed(22'h100000);
  assign T17894 = $signed(31'h4b730e70) * $signed(16'h1);
  assign T17895 = T10817[1'h0:1'h0];
  assign T17896 = T17905 ? twiddle4_2_415_real : twiddle4_2_414_real;
  assign twiddle4_2_414_real = T17899 + T17897;
  assign T17897 = $signed(T17898) / $signed(22'h100000);
  assign T17898 = $signed(31'h2434f332) * $signed(16'h0);
  assign T17899 = $signed(T17900) / $signed(22'h100000);
  assign T17900 = $signed(31'h4b39edca) * $signed(16'h1);
  assign twiddle4_2_415_real = T17903 + T17901;
  assign T17901 = $signed(T17902) / $signed(22'h100000);
  assign T17902 = $signed(31'h23e1e117) * $signed(16'h0);
  assign T17903 = $signed(T17904) / $signed(22'h100000);
  assign T17904 = $signed(31'h4b014f5b) * $signed(16'h1);
  assign T17905 = T10817[1'h0:1'h0];
  assign T17906 = T10817[1'h1:1'h1];
  assign T17907 = T10817[2'h2:2'h2];
  assign T17908 = T10817[2'h3:2'h3];
  assign T17909 = T10817[3'h4:3'h4];
  assign T17910 = T18141 ? T18015 : T17911;
  assign T17911 = T18014 ? T17958 : T17912;
  assign T17912 = T17957 ? T17935 : T17913;
  assign T17913 = T17934 ? T17924 : T17914;
  assign T17914 = T17923 ? twiddle4_2_417_real : twiddle4_2_416_real;
  assign twiddle4_2_416_real = T17917 + T17915;
  assign T17915 = $signed(T17916) / $signed(22'h100000);
  assign T17916 = $signed(31'h238e7673) * $signed(16'h0);
  assign T17917 = $signed(T17918) / $signed(22'h100000);
  assign T17918 = $signed(31'h4ac933ae) * $signed(16'h1);
  assign twiddle4_2_417_real = T17921 + T17919;
  assign T17919 = $signed(T17920) / $signed(22'h100000);
  assign T17920 = $signed(31'h233ab413) * $signed(16'h0);
  assign T17921 = $signed(T17922) / $signed(22'h100000);
  assign T17922 = $signed(31'h4a919b4e) * $signed(16'h1);
  assign T17923 = T10817[1'h0:1'h0];
  assign T17924 = T17933 ? twiddle4_2_419_real : twiddle4_2_418_real;
  assign twiddle4_2_418_real = T17927 + T17925;
  assign T17925 = $signed(T17926) / $signed(22'h100000);
  assign T17926 = $signed(31'h22e69ac7) * $signed(16'h0);
  assign T17927 = $signed(T17928) / $signed(22'h100000);
  assign T17928 = $signed(31'h4a5a86c4) * $signed(16'h1);
  assign twiddle4_2_419_real = T17931 + T17929;
  assign T17929 = $signed(T17930) / $signed(22'h100000);
  assign T17930 = $signed(31'h22922b5e) * $signed(16'h0);
  assign T17931 = $signed(T17932) / $signed(22'h100000);
  assign T17932 = $signed(31'h4a23f698) * $signed(16'h1);
  assign T17933 = T10817[1'h0:1'h0];
  assign T17934 = T10817[1'h1:1'h1];
  assign T17935 = T17956 ? T17946 : T17936;
  assign T17936 = T17945 ? twiddle4_2_421_real : twiddle4_2_420_real;
  assign twiddle4_2_420_real = T17939 + T17937;
  assign T17937 = $signed(T17938) / $signed(22'h100000);
  assign T17938 = $signed(31'h223d66a8) * $signed(16'h0);
  assign T17939 = $signed(T17940) / $signed(22'h100000);
  assign T17940 = $signed(31'h49edeb50) * $signed(16'h1);
  assign twiddle4_2_421_real = T17943 + T17941;
  assign T17941 = $signed(T17942) / $signed(22'h100000);
  assign T17942 = $signed(31'h21e84d76) * $signed(16'h0);
  assign T17943 = $signed(T17944) / $signed(22'h100000);
  assign T17944 = $signed(31'h49b86572) * $signed(16'h1);
  assign T17945 = T10817[1'h0:1'h0];
  assign T17946 = T17955 ? twiddle4_2_423_real : twiddle4_2_422_real;
  assign twiddle4_2_422_real = T17949 + T17947;
  assign T17947 = $signed(T17948) / $signed(22'h100000);
  assign T17948 = $signed(31'h2192e09a) * $signed(16'h0);
  assign T17949 = $signed(T17950) / $signed(22'h100000);
  assign T17950 = $signed(31'h49836583) * $signed(16'h1);
  assign twiddle4_2_423_real = T17953 + T17951;
  assign T17951 = $signed(T17952) / $signed(22'h100000);
  assign T17952 = $signed(31'h213d20e8) * $signed(16'h0);
  assign T17953 = $signed(T17954) / $signed(22'h100000);
  assign T17954 = $signed(31'h494eec03) * $signed(16'h1);
  assign T17955 = T10817[1'h0:1'h0];
  assign T17956 = T10817[1'h1:1'h1];
  assign T17957 = T10817[2'h2:2'h2];
  assign T17958 = T18013 ? T17983 : T17959;
  assign T17959 = T17982 ? T17970 : T17960;
  assign T17960 = T17969 ? twiddle4_2_425_real : twiddle4_2_424_real;
  assign twiddle4_2_424_real = T17963 + T17961;
  assign T17961 = $signed(T17962) / $signed(22'h100000);
  assign T17962 = $signed(31'h20e70f32) * $signed(16'h0);
  assign T17963 = $signed(T17964) / $signed(22'h100000);
  assign T17964 = $signed(31'h491af976) * $signed(16'h1);
  assign twiddle4_2_425_real = T17967 + T17965;
  assign T17965 = $signed(T17966) / $signed(22'h100000);
  assign T17966 = $signed(31'h2090ac4d) * $signed(16'h0);
  assign T17967 = $signed(T17968) / $signed(22'h100000);
  assign T17968 = $signed(31'h48e78e5c) * $signed(16'h1);
  assign T17969 = T10817[1'h0:1'h0];
  assign T17970 = T17981 ? twiddle4_2_427_real : twiddle4_2_426_real;
  assign twiddle4_2_426_real = T17973 + T17971;
  assign T17971 = $signed(T17972) / $signed(22'h100000);
  assign T17972 = $signed(31'h2039f90e) * $signed(16'h0);
  assign T17973 = $signed(T17974) / $signed(22'h100000);
  assign T17974 = $signed(31'h48b4ab32) * $signed(16'h1);
  assign twiddle4_2_427_real = T17979 + T17975;
  assign T17975 = {T17978, T17976};
  assign T17976 = $signed(T17977) / $signed(22'h100000);
  assign T17977 = $signed(30'h1fe2f64b) * $signed(16'h0);
  assign T17978 = T17976[6'h2d:6'h2d];
  assign T17979 = $signed(T17980) / $signed(22'h100000);
  assign T17980 = $signed(31'h48825077) * $signed(16'h1);
  assign T17981 = T10817[1'h0:1'h0];
  assign T17982 = T10817[1'h1:1'h1];
  assign T17983 = T18012 ? T17998 : T17984;
  assign T17984 = T17997 ? twiddle4_2_429_real : twiddle4_2_428_real;
  assign twiddle4_2_428_real = T17989 + T17985;
  assign T17985 = {T17988, T17986};
  assign T17986 = $signed(T17987) / $signed(22'h100000);
  assign T17987 = $signed(30'h1f8ba4db) * $signed(16'h0);
  assign T17988 = T17986[6'h2d:6'h2d];
  assign T17989 = $signed(T17990) / $signed(22'h100000);
  assign T17990 = $signed(31'h48507ea8) * $signed(16'h1);
  assign twiddle4_2_429_real = T17995 + T17991;
  assign T17991 = {T17994, T17992};
  assign T17992 = $signed(T17993) / $signed(22'h100000);
  assign T17993 = $signed(30'h1f340596) * $signed(16'h0);
  assign T17994 = T17992[6'h2d:6'h2d];
  assign T17995 = $signed(T17996) / $signed(22'h100000);
  assign T17996 = $signed(31'h481f363e) * $signed(16'h1);
  assign T17997 = T10817[1'h0:1'h0];
  assign T17998 = T18011 ? twiddle4_2_431_real : twiddle4_2_430_real;
  assign twiddle4_2_430_real = T18003 + T17999;
  assign T17999 = {T18002, T18000};
  assign T18000 = $signed(T18001) / $signed(22'h100000);
  assign T18001 = $signed(30'h1edc1952) * $signed(16'h0);
  assign T18002 = T18000[6'h2d:6'h2d];
  assign T18003 = $signed(T18004) / $signed(22'h100000);
  assign T18004 = $signed(31'h47ee77b4) * $signed(16'h1);
  assign twiddle4_2_431_real = T18009 + T18005;
  assign T18005 = {T18008, T18006};
  assign T18006 = $signed(T18007) / $signed(22'h100000);
  assign T18007 = $signed(30'h1e83e0ea) * $signed(16'h0);
  assign T18008 = T18006[6'h2d:6'h2d];
  assign T18009 = $signed(T18010) / $signed(22'h100000);
  assign T18010 = $signed(31'h47be4381) * $signed(16'h1);
  assign T18011 = T10817[1'h0:1'h0];
  assign T18012 = T10817[1'h1:1'h1];
  assign T18013 = T10817[2'h2:2'h2];
  assign T18014 = T10817[2'h3:2'h3];
  assign T18015 = T18140 ? T18078 : T18016;
  assign T18016 = T18077 ? T18047 : T18017;
  assign T18017 = T18046 ? T18032 : T18018;
  assign T18018 = T18031 ? twiddle4_2_433_real : twiddle4_2_432_real;
  assign twiddle4_2_432_real = T18023 + T18019;
  assign T18019 = {T18022, T18020};
  assign T18020 = $signed(T18021) / $signed(22'h100000);
  assign T18021 = $signed(30'h1e2b5d38) * $signed(16'h0);
  assign T18022 = T18020[6'h2d:6'h2d];
  assign T18023 = $signed(T18024) / $signed(22'h100000);
  assign T18024 = $signed(31'h478e9a1d) * $signed(16'h1);
  assign twiddle4_2_433_real = T18029 + T18025;
  assign T18025 = {T18028, T18026};
  assign T18026 = $signed(T18027) / $signed(22'h100000);
  assign T18027 = $signed(30'h1dd28f14) * $signed(16'h0);
  assign T18028 = T18026[6'h2d:6'h2d];
  assign T18029 = $signed(T18030) / $signed(22'h100000);
  assign T18030 = $signed(31'h475f7bfe) * $signed(16'h1);
  assign T18031 = T10817[1'h0:1'h0];
  assign T18032 = T18045 ? twiddle4_2_435_real : twiddle4_2_434_real;
  assign twiddle4_2_434_real = T18037 + T18033;
  assign T18033 = {T18036, T18034};
  assign T18034 = $signed(T18035) / $signed(22'h100000);
  assign T18035 = $signed(30'h1d79775b) * $signed(16'h0);
  assign T18036 = T18034[6'h2d:6'h2d];
  assign T18037 = $signed(T18038) / $signed(22'h100000);
  assign T18038 = $signed(31'h4730e997) * $signed(16'h1);
  assign twiddle4_2_435_real = T18043 + T18039;
  assign T18039 = {T18042, T18040};
  assign T18040 = $signed(T18041) / $signed(22'h100000);
  assign T18041 = $signed(30'h1d2016e8) * $signed(16'h0);
  assign T18042 = T18040[6'h2d:6'h2d];
  assign T18043 = $signed(T18044) / $signed(22'h100000);
  assign T18044 = $signed(31'h4702e35c) * $signed(16'h1);
  assign T18045 = T10817[1'h0:1'h0];
  assign T18046 = T10817[1'h1:1'h1];
  assign T18047 = T18076 ? T18062 : T18048;
  assign T18048 = T18061 ? twiddle4_2_437_real : twiddle4_2_436_real;
  assign twiddle4_2_436_real = T18053 + T18049;
  assign T18049 = {T18052, T18050};
  assign T18050 = $signed(T18051) / $signed(22'h100000);
  assign T18051 = $signed(30'h1cc66e99) * $signed(16'h0);
  assign T18052 = T18050[6'h2d:6'h2d];
  assign T18053 = $signed(T18054) / $signed(22'h100000);
  assign T18054 = $signed(31'h46d569be) * $signed(16'h1);
  assign twiddle4_2_437_real = T18059 + T18055;
  assign T18055 = {T18058, T18056};
  assign T18056 = $signed(T18057) / $signed(22'h100000);
  assign T18057 = $signed(30'h1c6c7f49) * $signed(16'h0);
  assign T18058 = T18056[6'h2d:6'h2d];
  assign T18059 = $signed(T18060) / $signed(22'h100000);
  assign T18060 = $signed(31'h46a87d2d) * $signed(16'h1);
  assign T18061 = T10817[1'h0:1'h0];
  assign T18062 = T18075 ? twiddle4_2_439_real : twiddle4_2_438_real;
  assign twiddle4_2_438_real = T18067 + T18063;
  assign T18063 = {T18066, T18064};
  assign T18064 = $signed(T18065) / $signed(22'h100000);
  assign T18065 = $signed(30'h1c1249d8) * $signed(16'h0);
  assign T18066 = T18064[6'h2d:6'h2d];
  assign T18067 = $signed(T18068) / $signed(22'h100000);
  assign T18068 = $signed(31'h467c1e19) * $signed(16'h1);
  assign twiddle4_2_439_real = T18073 + T18069;
  assign T18069 = {T18072, T18070};
  assign T18070 = $signed(T18071) / $signed(22'h100000);
  assign T18071 = $signed(30'h1bb7cf23) * $signed(16'h0);
  assign T18072 = T18070[6'h2d:6'h2d];
  assign T18073 = $signed(T18074) / $signed(22'h100000);
  assign T18074 = $signed(31'h46504ced) * $signed(16'h1);
  assign T18075 = T10817[1'h0:1'h0];
  assign T18076 = T10817[1'h1:1'h1];
  assign T18077 = T10817[2'h2:2'h2];
  assign T18078 = T18139 ? T18109 : T18079;
  assign T18079 = T18108 ? T18094 : T18080;
  assign T18080 = T18093 ? twiddle4_2_441_real : twiddle4_2_440_real;
  assign twiddle4_2_440_real = T18085 + T18081;
  assign T18081 = {T18084, T18082};
  assign T18082 = $signed(T18083) / $signed(22'h100000);
  assign T18083 = $signed(30'h1b5d1009) * $signed(16'h0);
  assign T18084 = T18082[6'h2d:6'h2d];
  assign T18085 = $signed(T18086) / $signed(22'h100000);
  assign T18086 = $signed(31'h46250a18) * $signed(16'h1);
  assign twiddle4_2_441_real = T18091 + T18087;
  assign T18087 = {T18090, T18088};
  assign T18088 = $signed(T18089) / $signed(22'h100000);
  assign T18089 = $signed(30'h1b020d6c) * $signed(16'h0);
  assign T18090 = T18088[6'h2d:6'h2d];
  assign T18091 = $signed(T18092) / $signed(22'h100000);
  assign T18092 = $signed(31'h45fa5603) * $signed(16'h1);
  assign T18093 = T10817[1'h0:1'h0];
  assign T18094 = T18107 ? twiddle4_2_443_real : twiddle4_2_442_real;
  assign twiddle4_2_442_real = T18099 + T18095;
  assign T18095 = {T18098, T18096};
  assign T18096 = $signed(T18097) / $signed(22'h100000);
  assign T18097 = $signed(30'h1aa6c82b) * $signed(16'h0);
  assign T18098 = T18096[6'h2d:6'h2d];
  assign T18099 = $signed(T18100) / $signed(22'h100000);
  assign T18100 = $signed(31'h45d03118) * $signed(16'h1);
  assign twiddle4_2_443_real = T18105 + T18101;
  assign T18101 = {T18104, T18102};
  assign T18102 = $signed(T18103) / $signed(22'h100000);
  assign T18103 = $signed(30'h1a4b4127) * $signed(16'h0);
  assign T18104 = T18102[6'h2d:6'h2d];
  assign T18105 = $signed(T18106) / $signed(22'h100000);
  assign T18106 = $signed(31'h45a69bbf) * $signed(16'h1);
  assign T18107 = T10817[1'h0:1'h0];
  assign T18108 = T10817[1'h1:1'h1];
  assign T18109 = T18138 ? T18124 : T18110;
  assign T18110 = T18123 ? twiddle4_2_445_real : twiddle4_2_444_real;
  assign twiddle4_2_444_real = T18115 + T18111;
  assign T18111 = {T18114, T18112};
  assign T18112 = $signed(T18113) / $signed(22'h100000);
  assign T18113 = $signed(30'h19ef7943) * $signed(16'h0);
  assign T18114 = T18112[6'h2d:6'h2d];
  assign T18115 = $signed(T18116) / $signed(22'h100000);
  assign T18116 = $signed(31'h457d965e) * $signed(16'h1);
  assign twiddle4_2_445_real = T18121 + T18117;
  assign T18117 = {T18120, T18118};
  assign T18118 = $signed(T18119) / $signed(22'h100000);
  assign T18119 = $signed(30'h19937161) * $signed(16'h0);
  assign T18120 = T18118[6'h2d:6'h2d];
  assign T18121 = $signed(T18122) / $signed(22'h100000);
  assign T18122 = $signed(31'h4555215b) * $signed(16'h1);
  assign T18123 = T10817[1'h0:1'h0];
  assign T18124 = T18137 ? twiddle4_2_447_real : twiddle4_2_446_real;
  assign twiddle4_2_446_real = T18129 + T18125;
  assign T18125 = {T18128, T18126};
  assign T18126 = $signed(T18127) / $signed(22'h100000);
  assign T18127 = $signed(30'h19372a63) * $signed(16'h0);
  assign T18128 = T18126[6'h2d:6'h2d];
  assign T18129 = $signed(T18130) / $signed(22'h100000);
  assign T18130 = $signed(31'h452d3d19) * $signed(16'h1);
  assign twiddle4_2_447_real = T18135 + T18131;
  assign T18131 = {T18134, T18132};
  assign T18132 = $signed(T18133) / $signed(22'h100000);
  assign T18133 = $signed(30'h18daa52e) * $signed(16'h0);
  assign T18134 = T18132[6'h2d:6'h2d];
  assign T18135 = $signed(T18136) / $signed(22'h100000);
  assign T18136 = $signed(31'h4505e9fb) * $signed(16'h1);
  assign T18137 = T10817[1'h0:1'h0];
  assign T18138 = T10817[1'h1:1'h1];
  assign T18139 = T10817[2'h2:2'h2];
  assign T18140 = T10817[2'h3:2'h3];
  assign T18141 = T10817[3'h4:3'h4];
  assign T18142 = T10817[3'h5:3'h5];
  assign T18143 = T18693 ? T18407 : T18144;
  assign T18144 = T18406 ? T18271 : T18145;
  assign T18145 = T18270 ? T18208 : T18146;
  assign T18146 = T18207 ? T18177 : T18147;
  assign T18147 = T18176 ? T18162 : T18148;
  assign T18148 = T18161 ? twiddle4_2_449_real : twiddle4_2_448_real;
  assign twiddle4_2_448_real = T18153 + T18149;
  assign T18149 = {T18152, T18150};
  assign T18150 = $signed(T18151) / $signed(22'h100000);
  assign T18151 = $signed(30'h187de2a6) * $signed(16'h0);
  assign T18152 = T18150[6'h2d:6'h2d];
  assign T18153 = $signed(T18154) / $signed(22'h100000);
  assign T18154 = $signed(31'h44df2862) * $signed(16'h1);
  assign twiddle4_2_449_real = T18159 + T18155;
  assign T18155 = {T18158, T18156};
  assign T18156 = $signed(T18157) / $signed(22'h100000);
  assign T18157 = $signed(30'h1820e3b0) * $signed(16'h0);
  assign T18158 = T18156[6'h2d:6'h2d];
  assign T18159 = $signed(T18160) / $signed(22'h100000);
  assign T18160 = $signed(31'h44b8f8ae) * $signed(16'h1);
  assign T18161 = T10817[1'h0:1'h0];
  assign T18162 = T18175 ? twiddle4_2_451_real : twiddle4_2_450_real;
  assign twiddle4_2_450_real = T18167 + T18163;
  assign T18163 = {T18166, T18164};
  assign T18164 = $signed(T18165) / $signed(22'h100000);
  assign T18165 = $signed(30'h17c3a931) * $signed(16'h0);
  assign T18166 = T18164[6'h2d:6'h2d];
  assign T18167 = $signed(T18168) / $signed(22'h100000);
  assign T18168 = $signed(31'h44935b3c) * $signed(16'h1);
  assign twiddle4_2_451_real = T18173 + T18169;
  assign T18169 = {T18172, T18170};
  assign T18170 = $signed(T18171) / $signed(22'h100000);
  assign T18171 = $signed(30'h1766340f) * $signed(16'h0);
  assign T18172 = T18170[6'h2d:6'h2d];
  assign T18173 = $signed(T18174) / $signed(22'h100000);
  assign T18174 = $signed(31'h446e506a) * $signed(16'h1);
  assign T18175 = T10817[1'h0:1'h0];
  assign T18176 = T10817[1'h1:1'h1];
  assign T18177 = T18206 ? T18192 : T18178;
  assign T18178 = T18191 ? twiddle4_2_453_real : twiddle4_2_452_real;
  assign twiddle4_2_452_real = T18183 + T18179;
  assign T18179 = {T18182, T18180};
  assign T18180 = $signed(T18181) / $signed(22'h100000);
  assign T18181 = $signed(30'h17088530) * $signed(16'h0);
  assign T18182 = T18180[6'h2d:6'h2d];
  assign T18183 = $signed(T18184) / $signed(22'h100000);
  assign T18184 = $signed(31'h4449d893) * $signed(16'h1);
  assign twiddle4_2_453_real = T18189 + T18185;
  assign T18185 = {T18188, T18186};
  assign T18186 = $signed(T18187) / $signed(22'h100000);
  assign T18187 = $signed(30'h16aa9d7d) * $signed(16'h0);
  assign T18188 = T18186[6'h2d:6'h2d];
  assign T18189 = $signed(T18190) / $signed(22'h100000);
  assign T18190 = $signed(31'h4425f411) * $signed(16'h1);
  assign T18191 = T10817[1'h0:1'h0];
  assign T18192 = T18205 ? twiddle4_2_455_real : twiddle4_2_454_real;
  assign twiddle4_2_454_real = T18197 + T18193;
  assign T18193 = {T18196, T18194};
  assign T18194 = $signed(T18195) / $signed(22'h100000);
  assign T18195 = $signed(30'h164c7ddd) * $signed(16'h0);
  assign T18196 = T18194[6'h2d:6'h2d];
  assign T18197 = $signed(T18198) / $signed(22'h100000);
  assign T18198 = $signed(31'h4402a33c) * $signed(16'h1);
  assign twiddle4_2_455_real = T18203 + T18199;
  assign T18199 = {T18202, T18200};
  assign T18200 = $signed(T18201) / $signed(22'h100000);
  assign T18201 = $signed(30'h15ee2737) * $signed(16'h0);
  assign T18202 = T18200[6'h2d:6'h2d];
  assign T18203 = $signed(T18204) / $signed(22'h100000);
  assign T18204 = $signed(31'h43dfe66c) * $signed(16'h1);
  assign T18205 = T10817[1'h0:1'h0];
  assign T18206 = T10817[1'h1:1'h1];
  assign T18207 = T10817[2'h2:2'h2];
  assign T18208 = T18269 ? T18239 : T18209;
  assign T18209 = T18238 ? T18224 : T18210;
  assign T18210 = T18223 ? twiddle4_2_457_real : twiddle4_2_456_real;
  assign twiddle4_2_456_real = T18215 + T18211;
  assign T18211 = {T18214, T18212};
  assign T18212 = $signed(T18213) / $signed(22'h100000);
  assign T18213 = $signed(30'h158f9a75) * $signed(16'h0);
  assign T18214 = T18212[6'h2d:6'h2d];
  assign T18215 = $signed(T18216) / $signed(22'h100000);
  assign T18216 = $signed(31'h43bdbdf7) * $signed(16'h1);
  assign twiddle4_2_457_real = T18221 + T18217;
  assign T18217 = {T18220, T18218};
  assign T18218 = $signed(T18219) / $signed(22'h100000);
  assign T18219 = $signed(30'h1530d880) * $signed(16'h0);
  assign T18220 = T18218[6'h2d:6'h2d];
  assign T18221 = $signed(T18222) / $signed(22'h100000);
  assign T18222 = $signed(31'h439c2a30) * $signed(16'h1);
  assign T18223 = T10817[1'h0:1'h0];
  assign T18224 = T18237 ? twiddle4_2_459_real : twiddle4_2_458_real;
  assign twiddle4_2_458_real = T18229 + T18225;
  assign T18225 = {T18228, T18226};
  assign T18226 = $signed(T18227) / $signed(22'h100000);
  assign T18227 = $signed(30'h14d1e242) * $signed(16'h0);
  assign T18228 = T18226[6'h2d:6'h2d];
  assign T18229 = $signed(T18230) / $signed(22'h100000);
  assign T18230 = $signed(31'h437b2b6a) * $signed(16'h1);
  assign twiddle4_2_459_real = T18235 + T18231;
  assign T18231 = {T18234, T18232};
  assign T18232 = $signed(T18233) / $signed(22'h100000);
  assign T18233 = $signed(30'h1472b8a5) * $signed(16'h0);
  assign T18234 = T18232[6'h2d:6'h2d];
  assign T18235 = $signed(T18236) / $signed(22'h100000);
  assign T18236 = $signed(31'h435ac1f8) * $signed(16'h1);
  assign T18237 = T10817[1'h0:1'h0];
  assign T18238 = T10817[1'h1:1'h1];
  assign T18239 = T18268 ? T18254 : T18240;
  assign T18240 = T18253 ? twiddle4_2_461_real : twiddle4_2_460_real;
  assign twiddle4_2_460_real = T18245 + T18241;
  assign T18241 = {T18244, T18242};
  assign T18242 = $signed(T18243) / $signed(22'h100000);
  assign T18243 = $signed(30'h14135c94) * $signed(16'h0);
  assign T18244 = T18242[6'h2d:6'h2d];
  assign T18245 = $signed(T18246) / $signed(22'h100000);
  assign T18246 = $signed(31'h433aee28) * $signed(16'h1);
  assign twiddle4_2_461_real = T18251 + T18247;
  assign T18247 = {T18250, T18248};
  assign T18248 = $signed(T18249) / $signed(22'h100000);
  assign T18249 = $signed(30'h13b3cefa) * $signed(16'h0);
  assign T18250 = T18248[6'h2d:6'h2d];
  assign T18251 = $signed(T18252) / $signed(22'h100000);
  assign T18252 = $signed(31'h431bb04a) * $signed(16'h1);
  assign T18253 = T10817[1'h0:1'h0];
  assign T18254 = T18267 ? twiddle4_2_463_real : twiddle4_2_462_real;
  assign twiddle4_2_462_real = T18259 + T18255;
  assign T18255 = {T18258, T18256};
  assign T18256 = $signed(T18257) / $signed(22'h100000);
  assign T18257 = $signed(30'h135410c2) * $signed(16'h0);
  assign T18258 = T18256[6'h2d:6'h2d];
  assign T18259 = $signed(T18260) / $signed(22'h100000);
  assign T18260 = $signed(31'h42fd08aa) * $signed(16'h1);
  assign twiddle4_2_463_real = T18265 + T18261;
  assign T18261 = {T18264, T18262};
  assign T18262 = $signed(T18263) / $signed(22'h100000);
  assign T18263 = $signed(30'h12f422da) * $signed(16'h0);
  assign T18264 = T18262[6'h2d:6'h2d];
  assign T18265 = $signed(T18266) / $signed(22'h100000);
  assign T18266 = $signed(31'h42def794) * $signed(16'h1);
  assign T18267 = T10817[1'h0:1'h0];
  assign T18268 = T10817[1'h1:1'h1];
  assign T18269 = T10817[2'h2:2'h2];
  assign T18270 = T10817[2'h3:2'h3];
  assign T18271 = T18405 ? T18335 : T18272;
  assign T18272 = T18334 ? T18303 : T18273;
  assign T18273 = T18302 ? T18288 : T18274;
  assign T18274 = T18287 ? twiddle4_2_465_real : twiddle4_2_464_real;
  assign twiddle4_2_464_real = T18279 + T18275;
  assign T18275 = {T18278, T18276};
  assign T18276 = $signed(T18277) / $signed(22'h100000);
  assign T18277 = $signed(30'h1294062e) * $signed(16'h0);
  assign T18278 = T18276[6'h2d:6'h2d];
  assign T18279 = $signed(T18280) / $signed(22'h100000);
  assign T18280 = $signed(31'h42c17d53) * $signed(16'h1);
  assign twiddle4_2_465_real = T18285 + T18281;
  assign T18281 = {T18284, T18282};
  assign T18282 = $signed(T18283) / $signed(22'h100000);
  assign T18283 = $signed(30'h1233bbab) * $signed(16'h0);
  assign T18284 = T18282[6'h2d:6'h2d];
  assign T18285 = $signed(T18286) / $signed(22'h100000);
  assign T18286 = $signed(31'h42a49a2f) * $signed(16'h1);
  assign T18287 = T10817[1'h0:1'h0];
  assign T18288 = T18301 ? twiddle4_2_467_real : twiddle4_2_466_real;
  assign twiddle4_2_466_real = T18293 + T18289;
  assign T18289 = {T18292, T18290};
  assign T18290 = $signed(T18291) / $signed(22'h100000);
  assign T18291 = $signed(30'h11d3443f) * $signed(16'h0);
  assign T18292 = T18290[6'h2d:6'h2d];
  assign T18293 = $signed(T18294) / $signed(22'h100000);
  assign T18294 = $signed(31'h42884e6f) * $signed(16'h1);
  assign twiddle4_2_467_real = T18299 + T18295;
  assign T18295 = {T18298, T18296};
  assign T18296 = $signed(T18297) / $signed(22'h100000);
  assign T18297 = $signed(30'h1172a0d7) * $signed(16'h0);
  assign T18298 = T18296[6'h2d:6'h2d];
  assign T18299 = $signed(T18300) / $signed(22'h100000);
  assign T18300 = $signed(31'h426c9a59) * $signed(16'h1);
  assign T18301 = T10817[1'h0:1'h0];
  assign T18302 = T10817[1'h1:1'h1];
  assign T18303 = T18333 ? T18318 : T18304;
  assign T18304 = T18317 ? twiddle4_2_469_real : twiddle4_2_468_real;
  assign twiddle4_2_468_real = T18309 + T18305;
  assign T18305 = {T18308, T18306};
  assign T18306 = $signed(T18307) / $signed(22'h100000);
  assign T18307 = $signed(30'h1111d262) * $signed(16'h0);
  assign T18308 = T18306[6'h2d:6'h2d];
  assign T18309 = $signed(T18310) / $signed(22'h100000);
  assign T18310 = $signed(31'h42517e32) * $signed(16'h1);
  assign twiddle4_2_469_real = T18315 + T18311;
  assign T18311 = {T18314, T18312};
  assign T18312 = $signed(T18313) / $signed(22'h100000);
  assign T18313 = $signed(30'h10b0d9cf) * $signed(16'h0);
  assign T18314 = T18312[6'h2d:6'h2d];
  assign T18315 = $signed(T18316) / $signed(22'h100000);
  assign T18316 = $signed(31'h4236fa3c) * $signed(16'h1);
  assign T18317 = T10817[1'h0:1'h0];
  assign T18318 = T18332 ? twiddle4_2_471_real : twiddle4_2_470_real;
  assign twiddle4_2_470_real = T18323 + T18319;
  assign T18319 = {T18322, T18320};
  assign T18320 = $signed(T18321) / $signed(22'h100000);
  assign T18321 = $signed(30'h104fb80e) * $signed(16'h0);
  assign T18322 = T18320[6'h2d:6'h2d];
  assign T18323 = $signed(T18324) / $signed(22'h100000);
  assign T18324 = $signed(31'h421d0eb9) * $signed(16'h1);
  assign twiddle4_2_471_real = T18330 + T18325;
  assign T18325 = {T18328, T18326};
  assign T18326 = $signed(T18327) / $signed(22'h100000);
  assign T18327 = $signed(29'hfee6e0d) * $signed(16'h0);
  assign T18328 = T18329 ? 2'h3 : 2'h0;
  assign T18329 = T18326[6'h2c:6'h2c];
  assign T18330 = $signed(T18331) / $signed(22'h100000);
  assign T18331 = $signed(31'h4203bbe8) * $signed(16'h1);
  assign T18332 = T10817[1'h0:1'h0];
  assign T18333 = T10817[1'h1:1'h1];
  assign T18334 = T10817[2'h2:2'h2];
  assign T18335 = T18404 ? T18370 : T18336;
  assign T18336 = T18369 ? T18353 : T18337;
  assign T18337 = T18352 ? twiddle4_2_473_real : twiddle4_2_472_real;
  assign twiddle4_2_472_real = T18343 + T18338;
  assign T18338 = {T18341, T18339};
  assign T18339 = $signed(T18340) / $signed(22'h100000);
  assign T18340 = $signed(29'hf8cfcbd) * $signed(16'h0);
  assign T18341 = T18342 ? 2'h3 : 2'h0;
  assign T18342 = T18339[6'h2c:6'h2c];
  assign T18343 = $signed(T18344) / $signed(22'h100000);
  assign T18344 = $signed(31'h41eb0209) * $signed(16'h1);
  assign twiddle4_2_473_real = T18350 + T18345;
  assign T18345 = {T18348, T18346};
  assign T18346 = $signed(T18347) / $signed(22'h100000);
  assign T18347 = $signed(29'hf2b650f) * $signed(16'h0);
  assign T18348 = T18349 ? 2'h3 : 2'h0;
  assign T18349 = T18346[6'h2c:6'h2c];
  assign T18350 = $signed(T18351) / $signed(22'h100000);
  assign T18351 = $signed(31'h41d2e159) * $signed(16'h1);
  assign T18352 = T10817[1'h0:1'h0];
  assign T18353 = T18368 ? twiddle4_2_475_real : twiddle4_2_474_real;
  assign twiddle4_2_474_real = T18359 + T18354;
  assign T18354 = {T18357, T18355};
  assign T18355 = $signed(T18356) / $signed(22'h100000);
  assign T18356 = $signed(29'hec9a7f2) * $signed(16'h0);
  assign T18357 = T18358 ? 2'h3 : 2'h0;
  assign T18358 = T18355[6'h2c:6'h2c];
  assign T18359 = $signed(T18360) / $signed(22'h100000);
  assign T18360 = $signed(31'h41bb5a12) * $signed(16'h1);
  assign twiddle4_2_475_real = T18366 + T18361;
  assign T18361 = {T18364, T18362};
  assign T18362 = $signed(T18363) / $signed(22'h100000);
  assign T18363 = $signed(29'he67c659) * $signed(16'h0);
  assign T18364 = T18365 ? 2'h3 : 2'h0;
  assign T18365 = T18362[6'h2c:6'h2c];
  assign T18366 = $signed(T18367) / $signed(22'h100000);
  assign T18367 = $signed(31'h41a46c6e) * $signed(16'h1);
  assign T18368 = T10817[1'h0:1'h0];
  assign T18369 = T10817[1'h1:1'h1];
  assign T18370 = T18403 ? T18387 : T18371;
  assign T18371 = T18386 ? twiddle4_2_477_real : twiddle4_2_476_real;
  assign twiddle4_2_476_real = T18377 + T18372;
  assign T18372 = {T18375, T18373};
  assign T18373 = $signed(T18374) / $signed(22'h100000);
  assign T18374 = $signed(29'he05c135) * $signed(16'h0);
  assign T18375 = T18376 ? 2'h3 : 2'h0;
  assign T18376 = T18373[6'h2c:6'h2c];
  assign T18377 = $signed(T18378) / $signed(22'h100000);
  assign T18378 = $signed(31'h418e18a8) * $signed(16'h1);
  assign twiddle4_2_477_real = T18384 + T18379;
  assign T18379 = {T18382, T18380};
  assign T18380 = $signed(T18381) / $signed(22'h100000);
  assign T18381 = $signed(29'hda39977) * $signed(16'h0);
  assign T18382 = T18383 ? 2'h3 : 2'h0;
  assign T18383 = T18380[6'h2c:6'h2c];
  assign T18384 = $signed(T18385) / $signed(22'h100000);
  assign T18385 = $signed(31'h41785ef5) * $signed(16'h1);
  assign T18386 = T10817[1'h0:1'h0];
  assign T18387 = T18402 ? twiddle4_2_479_real : twiddle4_2_478_real;
  assign twiddle4_2_478_real = T18393 + T18388;
  assign T18388 = {T18391, T18389};
  assign T18389 = $signed(T18390) / $signed(22'h100000);
  assign T18390 = $signed(29'hd415012) * $signed(16'h0);
  assign T18391 = T18392 ? 2'h3 : 2'h0;
  assign T18392 = T18389[6'h2c:6'h2c];
  assign T18393 = $signed(T18394) / $signed(22'h100000);
  assign T18394 = $signed(31'h41633f8a) * $signed(16'h1);
  assign twiddle4_2_479_real = T18400 + T18395;
  assign T18395 = {T18398, T18396};
  assign T18396 = $signed(T18397) / $signed(22'h100000);
  assign T18397 = $signed(29'hcdee5f9) * $signed(16'h0);
  assign T18398 = T18399 ? 2'h3 : 2'h0;
  assign T18399 = T18396[6'h2c:6'h2c];
  assign T18400 = $signed(T18401) / $signed(22'h100000);
  assign T18401 = $signed(31'h414eba9e) * $signed(16'h1);
  assign T18402 = T10817[1'h0:1'h0];
  assign T18403 = T10817[1'h1:1'h1];
  assign T18404 = T10817[2'h2:2'h2];
  assign T18405 = T10817[2'h3:2'h3];
  assign T18406 = T10817[3'h4:3'h4];
  assign T18407 = T18692 ? T18550 : T18408;
  assign T18408 = T18549 ? T18479 : T18409;
  assign T18409 = T18478 ? T18444 : T18410;
  assign T18410 = T18443 ? T18427 : T18411;
  assign T18411 = T18426 ? twiddle4_2_481_real : twiddle4_2_480_real;
  assign twiddle4_2_480_real = T18417 + T18412;
  assign T18412 = {T18415, T18413};
  assign T18413 = $signed(T18414) / $signed(22'h100000);
  assign T18414 = $signed(29'hc7c5c1e) * $signed(16'h0);
  assign T18415 = T18416 ? 2'h3 : 2'h0;
  assign T18416 = T18413[6'h2c:6'h2c];
  assign T18417 = $signed(T18418) / $signed(22'h100000);
  assign T18418 = $signed(31'h413ad061) * $signed(16'h1);
  assign twiddle4_2_481_real = T18424 + T18419;
  assign T18419 = {T18422, T18420};
  assign T18420 = $signed(T18421) / $signed(22'h100000);
  assign T18421 = $signed(29'hc19b374) * $signed(16'h0);
  assign T18422 = T18423 ? 2'h3 : 2'h0;
  assign T18423 = T18420[6'h2c:6'h2c];
  assign T18424 = $signed(T18425) / $signed(22'h100000);
  assign T18425 = $signed(31'h41278105) * $signed(16'h1);
  assign T18426 = T10817[1'h0:1'h0];
  assign T18427 = T18442 ? twiddle4_2_483_real : twiddle4_2_482_real;
  assign twiddle4_2_482_real = T18433 + T18428;
  assign T18428 = {T18431, T18429};
  assign T18429 = $signed(T18430) / $signed(22'h100000);
  assign T18430 = $signed(29'hbb6ecef) * $signed(16'h0);
  assign T18431 = T18432 ? 2'h3 : 2'h0;
  assign T18432 = T18429[6'h2c:6'h2c];
  assign T18433 = $signed(T18434) / $signed(22'h100000);
  assign T18434 = $signed(31'h4114ccb9) * $signed(16'h1);
  assign twiddle4_2_483_real = T18440 + T18435;
  assign T18435 = {T18438, T18436};
  assign T18436 = $signed(T18437) / $signed(22'h100000);
  assign T18437 = $signed(29'hb540982) * $signed(16'h0);
  assign T18438 = T18439 ? 2'h3 : 2'h0;
  assign T18439 = T18436[6'h2c:6'h2c];
  assign T18440 = $signed(T18441) / $signed(22'h100000);
  assign T18441 = $signed(31'h4102b3ad) * $signed(16'h1);
  assign T18442 = T10817[1'h0:1'h0];
  assign T18443 = T10817[1'h1:1'h1];
  assign T18444 = T18477 ? T18461 : T18445;
  assign T18445 = T18460 ? twiddle4_2_485_real : twiddle4_2_484_real;
  assign twiddle4_2_484_real = T18451 + T18446;
  assign T18446 = {T18449, T18447};
  assign T18447 = $signed(T18448) / $signed(22'h100000);
  assign T18448 = $signed(29'haf10a22) * $signed(16'h0);
  assign T18449 = T18450 ? 2'h3 : 2'h0;
  assign T18450 = T18447[6'h2c:6'h2c];
  assign T18451 = $signed(T18452) / $signed(22'h100000);
  assign T18452 = $signed(31'h40f1360c) * $signed(16'h1);
  assign twiddle4_2_485_real = T18458 + T18453;
  assign T18453 = {T18456, T18454};
  assign T18454 = $signed(T18455) / $signed(22'h100000);
  assign T18455 = $signed(29'ha8defc2) * $signed(16'h0);
  assign T18456 = T18457 ? 2'h3 : 2'h0;
  assign T18457 = T18454[6'h2c:6'h2c];
  assign T18458 = $signed(T18459) / $signed(22'h100000);
  assign T18459 = $signed(31'h40e05401) * $signed(16'h1);
  assign T18460 = T10817[1'h0:1'h0];
  assign T18461 = T18476 ? twiddle4_2_487_real : twiddle4_2_486_real;
  assign twiddle4_2_486_real = T18467 + T18462;
  assign T18462 = {T18465, T18463};
  assign T18463 = $signed(T18464) / $signed(22'h100000);
  assign T18464 = $signed(29'ha2abb58) * $signed(16'h0);
  assign T18465 = T18466 ? 2'h3 : 2'h0;
  assign T18466 = T18463[6'h2c:6'h2c];
  assign T18467 = $signed(T18468) / $signed(22'h100000);
  assign T18468 = $signed(31'h40d00db7) * $signed(16'h1);
  assign twiddle4_2_487_real = T18474 + T18469;
  assign T18469 = {T18472, T18470};
  assign T18470 = $signed(T18471) / $signed(22'h100000);
  assign T18471 = $signed(29'h9c76dd8) * $signed(16'h0);
  assign T18472 = T18473 ? 2'h3 : 2'h0;
  assign T18473 = T18470[6'h2c:6'h2c];
  assign T18474 = $signed(T18475) / $signed(22'h100000);
  assign T18475 = $signed(31'h40c06355) * $signed(16'h1);
  assign T18476 = T10817[1'h0:1'h0];
  assign T18477 = T10817[1'h1:1'h1];
  assign T18478 = T10817[2'h2:2'h2];
  assign T18479 = T18548 ? T18514 : T18480;
  assign T18480 = T18513 ? T18497 : T18481;
  assign T18481 = T18496 ? twiddle4_2_489_real : twiddle4_2_488_real;
  assign twiddle4_2_488_real = T18487 + T18482;
  assign T18482 = {T18485, T18483};
  assign T18483 = $signed(T18484) / $signed(22'h100000);
  assign T18484 = $signed(29'h9640837) * $signed(16'h0);
  assign T18485 = T18486 ? 2'h3 : 2'h0;
  assign T18486 = T18483[6'h2c:6'h2c];
  assign T18487 = $signed(T18488) / $signed(22'h100000);
  assign T18488 = $signed(31'h40b15502) * $signed(16'h1);
  assign twiddle4_2_489_real = T18494 + T18489;
  assign T18489 = {T18492, T18490};
  assign T18490 = $signed(T18491) / $signed(22'h100000);
  assign T18491 = $signed(29'h9008b6a) * $signed(16'h0);
  assign T18492 = T18493 ? 2'h3 : 2'h0;
  assign T18493 = T18490[6'h2c:6'h2c];
  assign T18494 = $signed(T18495) / $signed(22'h100000);
  assign T18495 = $signed(31'h40a2e2e4) * $signed(16'h1);
  assign T18496 = T10817[1'h0:1'h0];
  assign T18497 = T18512 ? twiddle4_2_491_real : twiddle4_2_490_real;
  assign twiddle4_2_490_real = T18503 + T18498;
  assign T18498 = {T18501, T18499};
  assign T18499 = $signed(T18500) / $signed(22'h100000);
  assign T18500 = $signed(29'h89cf867) * $signed(16'h0);
  assign T18501 = T18502 ? 2'h3 : 2'h0;
  assign T18502 = T18499[6'h2c:6'h2c];
  assign T18503 = $signed(T18504) / $signed(22'h100000);
  assign T18504 = $signed(31'h40950d1d) * $signed(16'h1);
  assign twiddle4_2_491_real = T18510 + T18505;
  assign T18505 = {T18508, T18506};
  assign T18506 = $signed(T18507) / $signed(22'h100000);
  assign T18507 = $signed(29'h8395023) * $signed(16'h0);
  assign T18508 = T18509 ? 2'h3 : 2'h0;
  assign T18509 = T18506[6'h2c:6'h2c];
  assign T18510 = $signed(T18511) / $signed(22'h100000);
  assign T18511 = $signed(31'h4087d3d1) * $signed(16'h1);
  assign T18512 = T10817[1'h0:1'h0];
  assign T18513 = T10817[1'h1:1'h1];
  assign T18514 = T18547 ? T18531 : T18515;
  assign T18515 = T18530 ? twiddle4_2_493_real : twiddle4_2_492_real;
  assign twiddle4_2_492_real = T18521 + T18516;
  assign T18516 = {T18519, T18517};
  assign T18517 = $signed(T18518) / $signed(22'h100000);
  assign T18518 = $signed(28'h7d59395) * $signed(16'h0);
  assign T18519 = T18520 ? 3'h7 : 3'h0;
  assign T18520 = T18517[6'h2b:6'h2b];
  assign T18521 = $signed(T18522) / $signed(22'h100000);
  assign T18522 = $signed(31'h407b371f) * $signed(16'h1);
  assign twiddle4_2_493_real = T18528 + T18523;
  assign T18523 = {T18526, T18524};
  assign T18524 = $signed(T18525) / $signed(22'h100000);
  assign T18525 = $signed(28'h771c3b2) * $signed(16'h0);
  assign T18526 = T18527 ? 3'h7 : 3'h0;
  assign T18527 = T18524[6'h2b:6'h2b];
  assign T18528 = $signed(T18529) / $signed(22'h100000);
  assign T18529 = $signed(31'h406f3727) * $signed(16'h1);
  assign T18530 = T10817[1'h0:1'h0];
  assign T18531 = T18546 ? twiddle4_2_495_real : twiddle4_2_494_real;
  assign twiddle4_2_494_real = T18537 + T18532;
  assign T18532 = {T18535, T18533};
  assign T18533 = $signed(T18534) / $signed(22'h100000);
  assign T18534 = $signed(28'h70de171) * $signed(16'h0);
  assign T18535 = T18536 ? 3'h7 : 3'h0;
  assign T18536 = T18533[6'h2b:6'h2b];
  assign T18537 = $signed(T18538) / $signed(22'h100000);
  assign T18538 = $signed(31'h4063d406) * $signed(16'h1);
  assign twiddle4_2_495_real = T18544 + T18539;
  assign T18539 = {T18542, T18540};
  assign T18540 = $signed(T18541) / $signed(22'h100000);
  assign T18541 = $signed(28'h6a9edc9) * $signed(16'h0);
  assign T18542 = T18543 ? 3'h7 : 3'h0;
  assign T18543 = T18540[6'h2b:6'h2b];
  assign T18544 = $signed(T18545) / $signed(22'h100000);
  assign T18545 = $signed(31'h40590dd8) * $signed(16'h1);
  assign T18546 = T10817[1'h0:1'h0];
  assign T18547 = T10817[1'h1:1'h1];
  assign T18548 = T10817[2'h2:2'h2];
  assign T18549 = T10817[2'h3:2'h3];
  assign T18550 = T18691 ? T18621 : T18551;
  assign T18551 = T18620 ? T18586 : T18552;
  assign T18552 = T18585 ? T18569 : T18553;
  assign T18553 = T18568 ? twiddle4_2_497_real : twiddle4_2_496_real;
  assign twiddle4_2_496_real = T18559 + T18554;
  assign T18554 = {T18557, T18555};
  assign T18555 = $signed(T18556) / $signed(22'h100000);
  assign T18556 = $signed(28'h645e9af) * $signed(16'h0);
  assign T18557 = T18558 ? 3'h7 : 3'h0;
  assign T18558 = T18555[6'h2b:6'h2b];
  assign T18559 = $signed(T18560) / $signed(22'h100000);
  assign T18560 = $signed(31'h404ee4b9) * $signed(16'h1);
  assign twiddle4_2_497_real = T18566 + T18561;
  assign T18561 = {T18564, T18562};
  assign T18562 = $signed(T18563) / $signed(22'h100000);
  assign T18563 = $signed(28'h5e1d61a) * $signed(16'h0);
  assign T18564 = T18565 ? 3'h7 : 3'h0;
  assign T18565 = T18562[6'h2b:6'h2b];
  assign T18566 = $signed(T18567) / $signed(22'h100000);
  assign T18567 = $signed(31'h404558c1) * $signed(16'h1);
  assign T18568 = T10817[1'h0:1'h0];
  assign T18569 = T18584 ? twiddle4_2_499_real : twiddle4_2_498_real;
  assign twiddle4_2_498_real = T18575 + T18570;
  assign T18570 = {T18573, T18571};
  assign T18571 = $signed(T18572) / $signed(22'h100000);
  assign T18572 = $signed(28'h57db402) * $signed(16'h0);
  assign T18573 = T18574 ? 3'h7 : 3'h0;
  assign T18574 = T18571[6'h2b:6'h2b];
  assign T18575 = $signed(T18576) / $signed(22'h100000);
  assign T18576 = $signed(31'h403c6a07) * $signed(16'h1);
  assign twiddle4_2_499_real = T18582 + T18577;
  assign T18577 = {T18580, T18578};
  assign T18578 = $signed(T18579) / $signed(22'h100000);
  assign T18579 = $signed(28'h519845e) * $signed(16'h0);
  assign T18580 = T18581 ? 3'h7 : 3'h0;
  assign T18581 = T18578[6'h2b:6'h2b];
  assign T18582 = $signed(T18583) / $signed(22'h100000);
  assign T18583 = $signed(31'h403418a2) * $signed(16'h1);
  assign T18584 = T10817[1'h0:1'h0];
  assign T18585 = T10817[1'h1:1'h1];
  assign T18586 = T18619 ? T18603 : T18587;
  assign T18587 = T18602 ? twiddle4_2_501_real : twiddle4_2_500_real;
  assign twiddle4_2_500_real = T18593 + T18588;
  assign T18588 = {T18591, T18589};
  assign T18589 = $signed(T18590) / $signed(22'h100000);
  assign T18590 = $signed(28'h4b54824) * $signed(16'h0);
  assign T18591 = T18592 ? 3'h7 : 3'h0;
  assign T18592 = T18589[6'h2b:6'h2b];
  assign T18593 = $signed(T18594) / $signed(22'h100000);
  assign T18594 = $signed(31'h402c64a6) * $signed(16'h1);
  assign twiddle4_2_501_real = T18600 + T18595;
  assign T18595 = {T18598, T18596};
  assign T18596 = $signed(T18597) / $signed(22'h100000);
  assign T18597 = $signed(28'h451004d) * $signed(16'h0);
  assign T18598 = T18599 ? 3'h7 : 3'h0;
  assign T18599 = T18596[6'h2b:6'h2b];
  assign T18600 = $signed(T18601) / $signed(22'h100000);
  assign T18601 = $signed(31'h40254e27) * $signed(16'h1);
  assign T18602 = T10817[1'h0:1'h0];
  assign T18603 = T18618 ? twiddle4_2_503_real : twiddle4_2_502_real;
  assign twiddle4_2_502_real = T18609 + T18604;
  assign T18604 = {T18607, T18605};
  assign T18605 = $signed(T18606) / $signed(22'h100000);
  assign T18606 = $signed(27'h3ecadcf) * $signed(16'h0);
  assign T18607 = T18608 ? 4'hf : 4'h0;
  assign T18608 = T18605[6'h2a:6'h2a];
  assign T18609 = $signed(T18610) / $signed(22'h100000);
  assign T18610 = $signed(31'h401ed535) * $signed(16'h1);
  assign twiddle4_2_503_real = T18616 + T18611;
  assign T18611 = {T18614, T18612};
  assign T18612 = $signed(T18613) / $signed(22'h100000);
  assign T18613 = $signed(27'h38851a2) * $signed(16'h0);
  assign T18614 = T18615 ? 4'hf : 4'h0;
  assign T18615 = T18612[6'h2a:6'h2a];
  assign T18616 = $signed(T18617) / $signed(22'h100000);
  assign T18617 = $signed(31'h4018f9e1) * $signed(16'h1);
  assign T18618 = T10817[1'h0:1'h0];
  assign T18619 = T10817[1'h1:1'h1];
  assign T18620 = T10817[2'h2:2'h2];
  assign T18621 = T18690 ? T18656 : T18622;
  assign T18622 = T18655 ? T18639 : T18623;
  assign T18623 = T18638 ? twiddle4_2_505_real : twiddle4_2_504_real;
  assign twiddle4_2_504_real = T18629 + T18624;
  assign T18624 = {T18627, T18625};
  assign T18625 = $signed(T18626) / $signed(22'h100000);
  assign T18626 = $signed(27'h323ecbe) * $signed(16'h0);
  assign T18627 = T18628 ? 4'hf : 4'h0;
  assign T18628 = T18625[6'h2a:6'h2a];
  assign T18629 = $signed(T18630) / $signed(22'h100000);
  assign T18630 = $signed(31'h4013bc3a) * $signed(16'h1);
  assign twiddle4_2_505_real = T18636 + T18631;
  assign T18631 = {T18634, T18632};
  assign T18632 = $signed(T18633) / $signed(22'h100000);
  assign T18633 = $signed(27'h2bf801a) * $signed(16'h0);
  assign T18634 = T18635 ? 4'hf : 4'h0;
  assign T18635 = T18632[6'h2a:6'h2a];
  assign T18636 = $signed(T18637) / $signed(22'h100000);
  assign T18637 = $signed(31'h400f1c4b) * $signed(16'h1);
  assign T18638 = T10817[1'h0:1'h0];
  assign T18639 = T18654 ? twiddle4_2_507_real : twiddle4_2_506_real;
  assign twiddle4_2_506_real = T18645 + T18640;
  assign T18640 = {T18643, T18641};
  assign T18641 = $signed(T18642) / $signed(22'h100000);
  assign T18642 = $signed(27'h25b0cae) * $signed(16'h0);
  assign T18643 = T18644 ? 4'hf : 4'h0;
  assign T18644 = T18641[6'h2a:6'h2a];
  assign T18645 = $signed(T18646) / $signed(22'h100000);
  assign T18646 = $signed(31'h400b1a21) * $signed(16'h1);
  assign twiddle4_2_507_real = T18652 + T18647;
  assign T18647 = {T18650, T18648};
  assign T18648 = $signed(T18649) / $signed(22'h100000);
  assign T18649 = $signed(26'h1f69373) * $signed(16'h0);
  assign T18650 = T18651 ? 5'h1f : 5'h0;
  assign T18651 = T18648[6'h29:6'h29];
  assign T18652 = $signed(T18653) / $signed(22'h100000);
  assign T18653 = $signed(31'h4007b5c5) * $signed(16'h1);
  assign T18654 = T10817[1'h0:1'h0];
  assign T18655 = T10817[1'h1:1'h1];
  assign T18656 = T18689 ? T18673 : T18657;
  assign T18657 = T18672 ? twiddle4_2_509_real : twiddle4_2_508_real;
  assign twiddle4_2_508_real = T18663 + T18658;
  assign T18658 = {T18661, T18659};
  assign T18659 = $signed(T18660) / $signed(22'h100000);
  assign T18660 = $signed(26'h192155f) * $signed(16'h0);
  assign T18661 = T18662 ? 5'h1f : 5'h0;
  assign T18662 = T18659[6'h29:6'h29];
  assign T18663 = $signed(T18664) / $signed(22'h100000);
  assign T18664 = $signed(31'h4004ef3f) * $signed(16'h1);
  assign twiddle4_2_509_real = T18670 + T18665;
  assign T18665 = {T18668, T18666};
  assign T18666 = $signed(T18667) / $signed(22'h100000);
  assign T18667 = $signed(26'h12d936b) * $signed(16'h0);
  assign T18668 = T18669 ? 5'h1f : 5'h0;
  assign T18669 = T18666[6'h29:6'h29];
  assign T18670 = $signed(T18671) / $signed(22'h100000);
  assign T18671 = $signed(31'h4002c698) * $signed(16'h1);
  assign T18672 = T10817[1'h0:1'h0];
  assign T18673 = T18688 ? twiddle4_2_511_real : twiddle4_2_510_real;
  assign twiddle4_2_510_real = T18679 + T18674;
  assign T18674 = {T18677, T18675};
  assign T18675 = $signed(T18676) / $signed(22'h100000);
  assign T18676 = $signed(25'hc90e8f) * $signed(16'h0);
  assign T18677 = T18678 ? 6'h3f : 6'h0;
  assign T18678 = T18675[6'h28:6'h28];
  assign T18679 = $signed(T18680) / $signed(22'h100000);
  assign T18680 = $signed(31'h40013bd3) * $signed(16'h1);
  assign twiddle4_2_511_real = T18686 + T18681;
  assign T18681 = {T18684, T18682};
  assign T18682 = $signed(T18683) / $signed(22'h100000);
  assign T18683 = $signed(24'h6487c3) * $signed(16'h0);
  assign T18684 = T18685 ? 7'h7f : 7'h0;
  assign T18685 = T18682[6'h27:6'h27];
  assign T18686 = $signed(T18687) / $signed(22'h100000);
  assign T18687 = $signed(31'h40004ef5) * $signed(16'h1);
  assign T18688 = T10817[1'h0:1'h0];
  assign T18689 = T10817[1'h1:1'h1];
  assign T18690 = T10817[2'h2:2'h2];
  assign T18691 = T10817[2'h3:2'h3];
  assign T18692 = T10817[3'h4:3'h4];
  assign T18693 = T10817[3'h5:3'h5];
  assign T18694 = T10817[3'h6:3'h6];
  assign T18695 = T17718[6'h2e:6'h2e];
  assign T18696 = T10817[3'h7:3'h7];
  assign T18697 = T10817[4'h8:4'h8];
  assign io_t4_1out_imag = T18698;
  assign T18698 = T18699[4'hf:1'h0];
  assign T18699 = T22635 ? T20677 : T18700;
  assign T18700 = T20676 ? T19822 : T18701;
  assign T18701 = T19821 ? T19290 : T18702;
  assign T18702 = T19289 ? T19001 : T18703;
  assign T18703 = T19000 ? T18856 : T18704;
  assign T18704 = T18855 ? T18783 : T18705;
  assign T18705 = T18782 ? T18746 : T18706;
  assign T18706 = T18745 ? T18727 : T18707;
  assign T18707 = T18724 ? T18715 : twiddle4_1_0_imag;
  assign twiddle4_1_0_imag = T18713 + T18708;
  assign T18708 = {T18711, T18709};
  assign T18709 = $signed(T18710) / $signed(22'h100000);
  assign T18710 = $signed(1'h0) * $signed(16'hffff);
  assign T18711 = T18712 ? 31'h7fffffff : 31'h0;
  assign T18712 = T18709[5'h10:5'h10];
  assign T18713 = $signed(T18714) / $signed(22'h100000);
  assign T18714 = $signed(32'h40000000) * $signed(16'h0);
  assign T18715 = {T18723, twiddle4_1_1_imag};
  assign twiddle4_1_1_imag = T18721 + T18716;
  assign T18716 = {T18719, T18717};
  assign T18717 = $signed(T18718) / $signed(22'h100000);
  assign T18718 = $signed(23'h3243f1) * $signed(16'hffff);
  assign T18719 = T18720 ? 8'hff : 8'h0;
  assign T18720 = T18717[6'h26:6'h26];
  assign T18721 = $signed(T18722) / $signed(22'h100000);
  assign T18722 = $signed(31'h3fffec42) * $signed(16'h0);
  assign T18723 = twiddle4_1_1_imag[6'h2e:6'h2e];
  assign T18724 = T18725[1'h0:1'h0];
  assign T18725 = T18726;
  assign T18726 = io_in4[4'h8:1'h0];
  assign T18727 = {T18744, T18728};
  assign T18728 = T18743 ? twiddle4_1_3_imag : twiddle4_1_2_imag;
  assign twiddle4_1_2_imag = T18734 + T18729;
  assign T18729 = {T18732, T18730};
  assign T18730 = $signed(T18731) / $signed(22'h100000);
  assign T18731 = $signed(24'h6487c3) * $signed(16'hffff);
  assign T18732 = T18733 ? 7'h7f : 7'h0;
  assign T18733 = T18730[6'h27:6'h27];
  assign T18734 = $signed(T18735) / $signed(22'h100000);
  assign T18735 = $signed(31'h3fffb10b) * $signed(16'h0);
  assign twiddle4_1_3_imag = T18741 + T18736;
  assign T18736 = {T18739, T18737};
  assign T18737 = $signed(T18738) / $signed(22'h100000);
  assign T18738 = $signed(25'h96cb58) * $signed(16'hffff);
  assign T18739 = T18740 ? 6'h3f : 6'h0;
  assign T18740 = T18737[6'h28:6'h28];
  assign T18741 = $signed(T18742) / $signed(22'h100000);
  assign T18742 = $signed(31'h3fff4e59) * $signed(16'h0);
  assign T18743 = T18725[1'h0:1'h0];
  assign T18744 = T18728[6'h2e:6'h2e];
  assign T18745 = T18725[1'h1:1'h1];
  assign T18746 = {T18781, T18747};
  assign T18747 = T18780 ? T18764 : T18748;
  assign T18748 = T18763 ? twiddle4_1_5_imag : twiddle4_1_4_imag;
  assign twiddle4_1_4_imag = T18754 + T18749;
  assign T18749 = {T18752, T18750};
  assign T18750 = $signed(T18751) / $signed(22'h100000);
  assign T18751 = $signed(25'hc90e8f) * $signed(16'hffff);
  assign T18752 = T18753 ? 6'h3f : 6'h0;
  assign T18753 = T18750[6'h28:6'h28];
  assign T18754 = $signed(T18755) / $signed(22'h100000);
  assign T18755 = $signed(31'h3ffec42d) * $signed(16'h0);
  assign twiddle4_1_5_imag = T18761 + T18756;
  assign T18756 = {T18759, T18757};
  assign T18757 = $signed(T18758) / $signed(22'h100000);
  assign T18758 = $signed(25'hfb514b) * $signed(16'hffff);
  assign T18759 = T18760 ? 6'h3f : 6'h0;
  assign T18760 = T18757[6'h28:6'h28];
  assign T18761 = $signed(T18762) / $signed(22'h100000);
  assign T18762 = $signed(31'h3ffe1287) * $signed(16'h0);
  assign T18763 = T18725[1'h0:1'h0];
  assign T18764 = T18779 ? twiddle4_1_7_imag : twiddle4_1_6_imag;
  assign twiddle4_1_6_imag = T18770 + T18765;
  assign T18765 = {T18768, T18766};
  assign T18766 = $signed(T18767) / $signed(22'h100000);
  assign T18767 = $signed(26'h12d936b) * $signed(16'hffff);
  assign T18768 = T18769 ? 5'h1f : 5'h0;
  assign T18769 = T18766[6'h29:6'h29];
  assign T18770 = $signed(T18771) / $signed(22'h100000);
  assign T18771 = $signed(31'h3ffd3968) * $signed(16'h0);
  assign twiddle4_1_7_imag = T18777 + T18772;
  assign T18772 = {T18775, T18773};
  assign T18773 = $signed(T18774) / $signed(22'h100000);
  assign T18774 = $signed(26'h15fd4d2) * $signed(16'hffff);
  assign T18775 = T18776 ? 5'h1f : 5'h0;
  assign T18776 = T18773[6'h29:6'h29];
  assign T18777 = $signed(T18778) / $signed(22'h100000);
  assign T18778 = $signed(31'h3ffc38d0) * $signed(16'h0);
  assign T18779 = T18725[1'h0:1'h0];
  assign T18780 = T18725[1'h1:1'h1];
  assign T18781 = T18747[6'h2e:6'h2e];
  assign T18782 = T18725[2'h2:2'h2];
  assign T18783 = {T18854, T18784};
  assign T18784 = T18853 ? T18819 : T18785;
  assign T18785 = T18818 ? T18802 : T18786;
  assign T18786 = T18801 ? twiddle4_1_9_imag : twiddle4_1_8_imag;
  assign twiddle4_1_8_imag = T18792 + T18787;
  assign T18787 = {T18790, T18788};
  assign T18788 = $signed(T18789) / $signed(22'h100000);
  assign T18789 = $signed(26'h192155f) * $signed(16'hffff);
  assign T18790 = T18791 ? 5'h1f : 5'h0;
  assign T18791 = T18788[6'h29:6'h29];
  assign T18792 = $signed(T18793) / $signed(22'h100000);
  assign T18793 = $signed(31'h3ffb10c1) * $signed(16'h0);
  assign twiddle4_1_9_imag = T18799 + T18794;
  assign T18794 = {T18797, T18795};
  assign T18795 = $signed(T18796) / $signed(22'h100000);
  assign T18796 = $signed(26'h1c454f4) * $signed(16'hffff);
  assign T18797 = T18798 ? 5'h1f : 5'h0;
  assign T18798 = T18795[6'h29:6'h29];
  assign T18799 = $signed(T18800) / $signed(22'h100000);
  assign T18800 = $signed(31'h3ff9c139) * $signed(16'h0);
  assign T18801 = T18725[1'h0:1'h0];
  assign T18802 = T18817 ? twiddle4_1_11_imag : twiddle4_1_10_imag;
  assign twiddle4_1_10_imag = T18808 + T18803;
  assign T18803 = {T18806, T18804};
  assign T18804 = $signed(T18805) / $signed(22'h100000);
  assign T18805 = $signed(26'h1f69373) * $signed(16'hffff);
  assign T18806 = T18807 ? 5'h1f : 5'h0;
  assign T18807 = T18804[6'h29:6'h29];
  assign T18808 = $signed(T18809) / $signed(22'h100000);
  assign T18809 = $signed(31'h3ff84a3b) * $signed(16'h0);
  assign twiddle4_1_11_imag = T18815 + T18810;
  assign T18810 = {T18813, T18811};
  assign T18811 = $signed(T18812) / $signed(22'h100000);
  assign T18812 = $signed(27'h228d0bb) * $signed(16'hffff);
  assign T18813 = T18814 ? 4'hf : 4'h0;
  assign T18814 = T18811[6'h2a:6'h2a];
  assign T18815 = $signed(T18816) / $signed(22'h100000);
  assign T18816 = $signed(31'h3ff6abc8) * $signed(16'h0);
  assign T18817 = T18725[1'h0:1'h0];
  assign T18818 = T18725[1'h1:1'h1];
  assign T18819 = T18852 ? T18836 : T18820;
  assign T18820 = T18835 ? twiddle4_1_13_imag : twiddle4_1_12_imag;
  assign twiddle4_1_12_imag = T18826 + T18821;
  assign T18821 = {T18824, T18822};
  assign T18822 = $signed(T18823) / $signed(22'h100000);
  assign T18823 = $signed(27'h25b0cae) * $signed(16'hffff);
  assign T18824 = T18825 ? 4'hf : 4'h0;
  assign T18825 = T18822[6'h2a:6'h2a];
  assign T18826 = $signed(T18827) / $signed(22'h100000);
  assign T18827 = $signed(31'h3ff4e5df) * $signed(16'h0);
  assign twiddle4_1_13_imag = T18833 + T18828;
  assign T18828 = {T18831, T18829};
  assign T18829 = $signed(T18830) / $signed(22'h100000);
  assign T18830 = $signed(27'h28d472d) * $signed(16'hffff);
  assign T18831 = T18832 ? 4'hf : 4'h0;
  assign T18832 = T18829[6'h2a:6'h2a];
  assign T18833 = $signed(T18834) / $signed(22'h100000);
  assign T18834 = $signed(31'h3ff2f884) * $signed(16'h0);
  assign T18835 = T18725[1'h0:1'h0];
  assign T18836 = T18851 ? twiddle4_1_15_imag : twiddle4_1_14_imag;
  assign twiddle4_1_14_imag = T18842 + T18837;
  assign T18837 = {T18840, T18838};
  assign T18838 = $signed(T18839) / $signed(22'h100000);
  assign T18839 = $signed(27'h2bf801a) * $signed(16'hffff);
  assign T18840 = T18841 ? 4'hf : 4'h0;
  assign T18841 = T18838[6'h2a:6'h2a];
  assign T18842 = $signed(T18843) / $signed(22'h100000);
  assign T18843 = $signed(31'h3ff0e3b5) * $signed(16'h0);
  assign twiddle4_1_15_imag = T18849 + T18844;
  assign T18844 = {T18847, T18845};
  assign T18845 = $signed(T18846) / $signed(22'h100000);
  assign T18846 = $signed(27'h2f1b754) * $signed(16'hffff);
  assign T18847 = T18848 ? 4'hf : 4'h0;
  assign T18848 = T18845[6'h2a:6'h2a];
  assign T18849 = $signed(T18850) / $signed(22'h100000);
  assign T18850 = $signed(31'h3feea776) * $signed(16'h0);
  assign T18851 = T18725[1'h0:1'h0];
  assign T18852 = T18725[1'h1:1'h1];
  assign T18853 = T18725[2'h2:2'h2];
  assign T18854 = T18784[6'h2e:6'h2e];
  assign T18855 = T18725[2'h3:2'h3];
  assign T18856 = {T18999, T18857};
  assign T18857 = T18998 ? T18928 : T18858;
  assign T18858 = T18927 ? T18893 : T18859;
  assign T18859 = T18892 ? T18876 : T18860;
  assign T18860 = T18875 ? twiddle4_1_17_imag : twiddle4_1_16_imag;
  assign twiddle4_1_16_imag = T18866 + T18861;
  assign T18861 = {T18864, T18862};
  assign T18862 = $signed(T18863) / $signed(22'h100000);
  assign T18863 = $signed(27'h323ecbe) * $signed(16'hffff);
  assign T18864 = T18865 ? 4'hf : 4'h0;
  assign T18865 = T18862[6'h2a:6'h2a];
  assign T18866 = $signed(T18867) / $signed(22'h100000);
  assign T18867 = $signed(31'h3fec43c6) * $signed(16'h0);
  assign twiddle4_1_17_imag = T18873 + T18868;
  assign T18868 = {T18871, T18869};
  assign T18869 = $signed(T18870) / $signed(22'h100000);
  assign T18870 = $signed(27'h3562037) * $signed(16'hffff);
  assign T18871 = T18872 ? 4'hf : 4'h0;
  assign T18872 = T18869[6'h2a:6'h2a];
  assign T18873 = $signed(T18874) / $signed(22'h100000);
  assign T18874 = $signed(31'h3fe9b8a9) * $signed(16'h0);
  assign T18875 = T18725[1'h0:1'h0];
  assign T18876 = T18891 ? twiddle4_1_19_imag : twiddle4_1_18_imag;
  assign twiddle4_1_18_imag = T18882 + T18877;
  assign T18877 = {T18880, T18878};
  assign T18878 = $signed(T18879) / $signed(22'h100000);
  assign T18879 = $signed(27'h38851a2) * $signed(16'hffff);
  assign T18880 = T18881 ? 4'hf : 4'h0;
  assign T18881 = T18878[6'h2a:6'h2a];
  assign T18882 = $signed(T18883) / $signed(22'h100000);
  assign T18883 = $signed(31'h3fe7061f) * $signed(16'h0);
  assign twiddle4_1_19_imag = T18889 + T18884;
  assign T18884 = {T18887, T18885};
  assign T18885 = $signed(T18886) / $signed(22'h100000);
  assign T18886 = $signed(27'h3ba80df) * $signed(16'hffff);
  assign T18887 = T18888 ? 4'hf : 4'h0;
  assign T18888 = T18885[6'h2a:6'h2a];
  assign T18889 = $signed(T18890) / $signed(22'h100000);
  assign T18890 = $signed(31'h3fe42c29) * $signed(16'h0);
  assign T18891 = T18725[1'h0:1'h0];
  assign T18892 = T18725[1'h1:1'h1];
  assign T18893 = T18926 ? T18910 : T18894;
  assign T18894 = T18909 ? twiddle4_1_21_imag : twiddle4_1_20_imag;
  assign twiddle4_1_20_imag = T18900 + T18895;
  assign T18895 = {T18898, T18896};
  assign T18896 = $signed(T18897) / $signed(22'h100000);
  assign T18897 = $signed(27'h3ecadcf) * $signed(16'hffff);
  assign T18898 = T18899 ? 4'hf : 4'h0;
  assign T18899 = T18896[6'h2a:6'h2a];
  assign T18900 = $signed(T18901) / $signed(22'h100000);
  assign T18901 = $signed(31'h3fe12acb) * $signed(16'h0);
  assign twiddle4_1_21_imag = T18907 + T18902;
  assign T18902 = {T18905, T18903};
  assign T18903 = $signed(T18904) / $signed(22'h100000);
  assign T18904 = $signed(28'h41ed853) * $signed(16'hffff);
  assign T18905 = T18906 ? 3'h7 : 3'h0;
  assign T18906 = T18903[6'h2b:6'h2b];
  assign T18907 = $signed(T18908) / $signed(22'h100000);
  assign T18908 = $signed(31'h3fde0205) * $signed(16'h0);
  assign T18909 = T18725[1'h0:1'h0];
  assign T18910 = T18925 ? twiddle4_1_23_imag : twiddle4_1_22_imag;
  assign twiddle4_1_22_imag = T18916 + T18911;
  assign T18911 = {T18914, T18912};
  assign T18912 = $signed(T18913) / $signed(22'h100000);
  assign T18913 = $signed(28'h451004d) * $signed(16'hffff);
  assign T18914 = T18915 ? 3'h7 : 3'h0;
  assign T18915 = T18912[6'h2b:6'h2b];
  assign T18916 = $signed(T18917) / $signed(22'h100000);
  assign T18917 = $signed(31'h3fdab1d9) * $signed(16'h0);
  assign twiddle4_1_23_imag = T18923 + T18918;
  assign T18918 = {T18921, T18919};
  assign T18919 = $signed(T18920) / $signed(22'h100000);
  assign T18920 = $signed(28'h483259d) * $signed(16'hffff);
  assign T18921 = T18922 ? 3'h7 : 3'h0;
  assign T18922 = T18919[6'h2b:6'h2b];
  assign T18923 = $signed(T18924) / $signed(22'h100000);
  assign T18924 = $signed(31'h3fd73a4a) * $signed(16'h0);
  assign T18925 = T18725[1'h0:1'h0];
  assign T18926 = T18725[1'h1:1'h1];
  assign T18927 = T18725[2'h2:2'h2];
  assign T18928 = T18997 ? T18963 : T18929;
  assign T18929 = T18962 ? T18946 : T18930;
  assign T18930 = T18945 ? twiddle4_1_25_imag : twiddle4_1_24_imag;
  assign twiddle4_1_24_imag = T18936 + T18931;
  assign T18931 = {T18934, T18932};
  assign T18932 = $signed(T18933) / $signed(22'h100000);
  assign T18933 = $signed(28'h4b54824) * $signed(16'hffff);
  assign T18934 = T18935 ? 3'h7 : 3'h0;
  assign T18935 = T18932[6'h2b:6'h2b];
  assign T18936 = $signed(T18937) / $signed(22'h100000);
  assign T18937 = $signed(31'h3fd39b5a) * $signed(16'h0);
  assign twiddle4_1_25_imag = T18943 + T18938;
  assign T18938 = {T18941, T18939};
  assign T18939 = $signed(T18940) / $signed(22'h100000);
  assign T18940 = $signed(28'h4e767c4) * $signed(16'hffff);
  assign T18941 = T18942 ? 3'h7 : 3'h0;
  assign T18942 = T18939[6'h2b:6'h2b];
  assign T18943 = $signed(T18944) / $signed(22'h100000);
  assign T18944 = $signed(31'h3fcfd50a) * $signed(16'h0);
  assign T18945 = T18725[1'h0:1'h0];
  assign T18946 = T18961 ? twiddle4_1_27_imag : twiddle4_1_26_imag;
  assign twiddle4_1_26_imag = T18952 + T18947;
  assign T18947 = {T18950, T18948};
  assign T18948 = $signed(T18949) / $signed(22'h100000);
  assign T18949 = $signed(28'h519845e) * $signed(16'hffff);
  assign T18950 = T18951 ? 3'h7 : 3'h0;
  assign T18951 = T18948[6'h2b:6'h2b];
  assign T18952 = $signed(T18953) / $signed(22'h100000);
  assign T18953 = $signed(31'h3fcbe75e) * $signed(16'h0);
  assign twiddle4_1_27_imag = T18959 + T18954;
  assign T18954 = {T18957, T18955};
  assign T18955 = $signed(T18956) / $signed(22'h100000);
  assign T18956 = $signed(28'h54b9dd2) * $signed(16'hffff);
  assign T18957 = T18958 ? 3'h7 : 3'h0;
  assign T18958 = T18955[6'h2b:6'h2b];
  assign T18959 = $signed(T18960) / $signed(22'h100000);
  assign T18960 = $signed(31'h3fc7d257) * $signed(16'h0);
  assign T18961 = T18725[1'h0:1'h0];
  assign T18962 = T18725[1'h1:1'h1];
  assign T18963 = T18996 ? T18980 : T18964;
  assign T18964 = T18979 ? twiddle4_1_29_imag : twiddle4_1_28_imag;
  assign twiddle4_1_28_imag = T18970 + T18965;
  assign T18965 = {T18968, T18966};
  assign T18966 = $signed(T18967) / $signed(22'h100000);
  assign T18967 = $signed(28'h57db402) * $signed(16'hffff);
  assign T18968 = T18969 ? 3'h7 : 3'h0;
  assign T18969 = T18966[6'h2b:6'h2b];
  assign T18970 = $signed(T18971) / $signed(22'h100000);
  assign T18971 = $signed(31'h3fc395f9) * $signed(16'h0);
  assign twiddle4_1_29_imag = T18977 + T18972;
  assign T18972 = {T18975, T18973};
  assign T18973 = $signed(T18974) / $signed(22'h100000);
  assign T18974 = $signed(28'h5afc6cf) * $signed(16'hffff);
  assign T18975 = T18976 ? 3'h7 : 3'h0;
  assign T18976 = T18973[6'h2b:6'h2b];
  assign T18977 = $signed(T18978) / $signed(22'h100000);
  assign T18978 = $signed(31'h3fbf3245) * $signed(16'h0);
  assign T18979 = T18725[1'h0:1'h0];
  assign T18980 = T18995 ? twiddle4_1_31_imag : twiddle4_1_30_imag;
  assign twiddle4_1_30_imag = T18986 + T18981;
  assign T18981 = {T18984, T18982};
  assign T18982 = $signed(T18983) / $signed(22'h100000);
  assign T18983 = $signed(28'h5e1d61a) * $signed(16'hffff);
  assign T18984 = T18985 ? 3'h7 : 3'h0;
  assign T18985 = T18982[6'h2b:6'h2b];
  assign T18986 = $signed(T18987) / $signed(22'h100000);
  assign T18987 = $signed(31'h3fbaa73f) * $signed(16'h0);
  assign twiddle4_1_31_imag = T18993 + T18988;
  assign T18988 = {T18991, T18989};
  assign T18989 = $signed(T18990) / $signed(22'h100000);
  assign T18990 = $signed(28'h613e1c4) * $signed(16'hffff);
  assign T18991 = T18992 ? 3'h7 : 3'h0;
  assign T18992 = T18989[6'h2b:6'h2b];
  assign T18993 = $signed(T18994) / $signed(22'h100000);
  assign T18994 = $signed(31'h3fb5f4ea) * $signed(16'h0);
  assign T18995 = T18725[1'h0:1'h0];
  assign T18996 = T18725[1'h1:1'h1];
  assign T18997 = T18725[2'h2:2'h2];
  assign T18998 = T18725[2'h3:2'h3];
  assign T18999 = T18857[6'h2e:6'h2e];
  assign T19000 = T18725[3'h4:3'h4];
  assign T19001 = {T19288, T19002};
  assign T19002 = T19287 ? T19145 : T19003;
  assign T19003 = T19144 ? T19074 : T19004;
  assign T19004 = T19073 ? T19039 : T19005;
  assign T19005 = T19038 ? T19022 : T19006;
  assign T19006 = T19021 ? twiddle4_1_33_imag : twiddle4_1_32_imag;
  assign twiddle4_1_32_imag = T19012 + T19007;
  assign T19007 = {T19010, T19008};
  assign T19008 = $signed(T19009) / $signed(22'h100000);
  assign T19009 = $signed(28'h645e9af) * $signed(16'hffff);
  assign T19010 = T19011 ? 3'h7 : 3'h0;
  assign T19011 = T19008[6'h2b:6'h2b];
  assign T19012 = $signed(T19013) / $signed(22'h100000);
  assign T19013 = $signed(31'h3fb11b47) * $signed(16'h0);
  assign twiddle4_1_33_imag = T19019 + T19014;
  assign T19014 = {T19017, T19015};
  assign T19015 = $signed(T19016) / $signed(22'h100000);
  assign T19016 = $signed(28'h677edba) * $signed(16'hffff);
  assign T19017 = T19018 ? 3'h7 : 3'h0;
  assign T19018 = T19015[6'h2b:6'h2b];
  assign T19019 = $signed(T19020) / $signed(22'h100000);
  assign T19020 = $signed(31'h3fac1a5b) * $signed(16'h0);
  assign T19021 = T18725[1'h0:1'h0];
  assign T19022 = T19037 ? twiddle4_1_35_imag : twiddle4_1_34_imag;
  assign twiddle4_1_34_imag = T19028 + T19023;
  assign T19023 = {T19026, T19024};
  assign T19024 = $signed(T19025) / $signed(22'h100000);
  assign T19025 = $signed(28'h6a9edc9) * $signed(16'hffff);
  assign T19026 = T19027 ? 3'h7 : 3'h0;
  assign T19027 = T19024[6'h2b:6'h2b];
  assign T19028 = $signed(T19029) / $signed(22'h100000);
  assign T19029 = $signed(31'h3fa6f228) * $signed(16'h0);
  assign twiddle4_1_35_imag = T19035 + T19030;
  assign T19030 = {T19033, T19031};
  assign T19031 = $signed(T19032) / $signed(22'h100000);
  assign T19032 = $signed(28'h6dbe9bb) * $signed(16'hffff);
  assign T19033 = T19034 ? 3'h7 : 3'h0;
  assign T19034 = T19031[6'h2b:6'h2b];
  assign T19035 = $signed(T19036) / $signed(22'h100000);
  assign T19036 = $signed(31'h3fa1a2b1) * $signed(16'h0);
  assign T19037 = T18725[1'h0:1'h0];
  assign T19038 = T18725[1'h1:1'h1];
  assign T19039 = T19072 ? T19056 : T19040;
  assign T19040 = T19055 ? twiddle4_1_37_imag : twiddle4_1_36_imag;
  assign twiddle4_1_36_imag = T19046 + T19041;
  assign T19041 = {T19044, T19042};
  assign T19042 = $signed(T19043) / $signed(22'h100000);
  assign T19043 = $signed(28'h70de171) * $signed(16'hffff);
  assign T19044 = T19045 ? 3'h7 : 3'h0;
  assign T19045 = T19042[6'h2b:6'h2b];
  assign T19046 = $signed(T19047) / $signed(22'h100000);
  assign T19047 = $signed(31'h3f9c2bfa) * $signed(16'h0);
  assign twiddle4_1_37_imag = T19053 + T19048;
  assign T19048 = {T19051, T19049};
  assign T19049 = $signed(T19050) / $signed(22'h100000);
  assign T19050 = $signed(28'h73fd4ce) * $signed(16'hffff);
  assign T19051 = T19052 ? 3'h7 : 3'h0;
  assign T19052 = T19049[6'h2b:6'h2b];
  assign T19053 = $signed(T19054) / $signed(22'h100000);
  assign T19054 = $signed(31'h3f968e07) * $signed(16'h0);
  assign T19055 = T18725[1'h0:1'h0];
  assign T19056 = T19071 ? twiddle4_1_39_imag : twiddle4_1_38_imag;
  assign twiddle4_1_38_imag = T19062 + T19057;
  assign T19057 = {T19060, T19058};
  assign T19058 = $signed(T19059) / $signed(22'h100000);
  assign T19059 = $signed(28'h771c3b2) * $signed(16'hffff);
  assign T19060 = T19061 ? 3'h7 : 3'h0;
  assign T19061 = T19058[6'h2b:6'h2b];
  assign T19062 = $signed(T19063) / $signed(22'h100000);
  assign T19063 = $signed(31'h3f90c8d9) * $signed(16'h0);
  assign twiddle4_1_39_imag = T19069 + T19064;
  assign T19064 = {T19067, T19065};
  assign T19065 = $signed(T19066) / $signed(22'h100000);
  assign T19066 = $signed(28'h7a3adff) * $signed(16'hffff);
  assign T19067 = T19068 ? 3'h7 : 3'h0;
  assign T19068 = T19065[6'h2b:6'h2b];
  assign T19069 = $signed(T19070) / $signed(22'h100000);
  assign T19070 = $signed(31'h3f8adc76) * $signed(16'h0);
  assign T19071 = T18725[1'h0:1'h0];
  assign T19072 = T18725[1'h1:1'h1];
  assign T19073 = T18725[2'h2:2'h2];
  assign T19074 = T19143 ? T19109 : T19075;
  assign T19075 = T19108 ? T19092 : T19076;
  assign T19076 = T19091 ? twiddle4_1_41_imag : twiddle4_1_40_imag;
  assign twiddle4_1_40_imag = T19082 + T19077;
  assign T19077 = {T19080, T19078};
  assign T19078 = $signed(T19079) / $signed(22'h100000);
  assign T19079 = $signed(28'h7d59395) * $signed(16'hffff);
  assign T19080 = T19081 ? 3'h7 : 3'h0;
  assign T19081 = T19078[6'h2b:6'h2b];
  assign T19082 = $signed(T19083) / $signed(22'h100000);
  assign T19083 = $signed(31'h3f84c8e1) * $signed(16'h0);
  assign twiddle4_1_41_imag = T19089 + T19084;
  assign T19084 = {T19087, T19085};
  assign T19085 = $signed(T19086) / $signed(22'h100000);
  assign T19086 = $signed(29'h8077456) * $signed(16'hffff);
  assign T19087 = T19088 ? 2'h3 : 2'h0;
  assign T19088 = T19085[6'h2c:6'h2c];
  assign T19089 = $signed(T19090) / $signed(22'h100000);
  assign T19090 = $signed(31'h3f7e8e1e) * $signed(16'h0);
  assign T19091 = T18725[1'h0:1'h0];
  assign T19092 = T19107 ? twiddle4_1_43_imag : twiddle4_1_42_imag;
  assign twiddle4_1_42_imag = T19098 + T19093;
  assign T19093 = {T19096, T19094};
  assign T19094 = $signed(T19095) / $signed(22'h100000);
  assign T19095 = $signed(29'h8395023) * $signed(16'hffff);
  assign T19096 = T19097 ? 2'h3 : 2'h0;
  assign T19097 = T19094[6'h2c:6'h2c];
  assign T19098 = $signed(T19099) / $signed(22'h100000);
  assign T19099 = $signed(31'h3f782c2f) * $signed(16'h0);
  assign twiddle4_1_43_imag = T19105 + T19100;
  assign T19100 = {T19103, T19101};
  assign T19101 = $signed(T19102) / $signed(22'h100000);
  assign T19102 = $signed(29'h86b26de) * $signed(16'hffff);
  assign T19103 = T19104 ? 2'h3 : 2'h0;
  assign T19104 = T19101[6'h2c:6'h2c];
  assign T19105 = $signed(T19106) / $signed(22'h100000);
  assign T19106 = $signed(31'h3f71a31a) * $signed(16'h0);
  assign T19107 = T18725[1'h0:1'h0];
  assign T19108 = T18725[1'h1:1'h1];
  assign T19109 = T19142 ? T19126 : T19110;
  assign T19110 = T19125 ? twiddle4_1_45_imag : twiddle4_1_44_imag;
  assign twiddle4_1_44_imag = T19116 + T19111;
  assign T19111 = {T19114, T19112};
  assign T19112 = $signed(T19113) / $signed(22'h100000);
  assign T19113 = $signed(29'h89cf867) * $signed(16'hffff);
  assign T19114 = T19115 ? 2'h3 : 2'h0;
  assign T19115 = T19112[6'h2c:6'h2c];
  assign T19116 = $signed(T19117) / $signed(22'h100000);
  assign T19117 = $signed(31'h3f6af2e3) * $signed(16'h0);
  assign twiddle4_1_45_imag = T19123 + T19118;
  assign T19118 = {T19121, T19119};
  assign T19119 = $signed(T19120) / $signed(22'h100000);
  assign T19120 = $signed(29'h8cec4a0) * $signed(16'hffff);
  assign T19121 = T19122 ? 2'h3 : 2'h0;
  assign T19122 = T19119[6'h2c:6'h2c];
  assign T19123 = $signed(T19124) / $signed(22'h100000);
  assign T19124 = $signed(31'h3f641b8d) * $signed(16'h0);
  assign T19125 = T18725[1'h0:1'h0];
  assign T19126 = T19141 ? twiddle4_1_47_imag : twiddle4_1_46_imag;
  assign twiddle4_1_46_imag = T19132 + T19127;
  assign T19127 = {T19130, T19128};
  assign T19128 = $signed(T19129) / $signed(22'h100000);
  assign T19129 = $signed(29'h9008b6a) * $signed(16'hffff);
  assign T19130 = T19131 ? 2'h3 : 2'h0;
  assign T19131 = T19128[6'h2c:6'h2c];
  assign T19132 = $signed(T19133) / $signed(22'h100000);
  assign T19133 = $signed(31'h3f5d1d1c) * $signed(16'h0);
  assign twiddle4_1_47_imag = T19139 + T19134;
  assign T19134 = {T19137, T19135};
  assign T19135 = $signed(T19136) / $signed(22'h100000);
  assign T19136 = $signed(29'h9324ca6) * $signed(16'hffff);
  assign T19137 = T19138 ? 2'h3 : 2'h0;
  assign T19138 = T19135[6'h2c:6'h2c];
  assign T19139 = $signed(T19140) / $signed(22'h100000);
  assign T19140 = $signed(31'h3f55f796) * $signed(16'h0);
  assign T19141 = T18725[1'h0:1'h0];
  assign T19142 = T18725[1'h1:1'h1];
  assign T19143 = T18725[2'h2:2'h2];
  assign T19144 = T18725[2'h3:2'h3];
  assign T19145 = T19286 ? T19216 : T19146;
  assign T19146 = T19215 ? T19181 : T19147;
  assign T19147 = T19180 ? T19164 : T19148;
  assign T19148 = T19163 ? twiddle4_1_49_imag : twiddle4_1_48_imag;
  assign twiddle4_1_48_imag = T19154 + T19149;
  assign T19149 = {T19152, T19150};
  assign T19150 = $signed(T19151) / $signed(22'h100000);
  assign T19151 = $signed(29'h9640837) * $signed(16'hffff);
  assign T19152 = T19153 ? 2'h3 : 2'h0;
  assign T19153 = T19150[6'h2c:6'h2c];
  assign T19154 = $signed(T19155) / $signed(22'h100000);
  assign T19155 = $signed(31'h3f4eaafe) * $signed(16'h0);
  assign twiddle4_1_49_imag = T19161 + T19156;
  assign T19156 = {T19159, T19157};
  assign T19157 = $signed(T19158) / $signed(22'h100000);
  assign T19158 = $signed(29'h995bdfc) * $signed(16'hffff);
  assign T19159 = T19160 ? 2'h3 : 2'h0;
  assign T19160 = T19157[6'h2c:6'h2c];
  assign T19161 = $signed(T19162) / $signed(22'h100000);
  assign T19162 = $signed(31'h3f473758) * $signed(16'h0);
  assign T19163 = T18725[1'h0:1'h0];
  assign T19164 = T19179 ? twiddle4_1_51_imag : twiddle4_1_50_imag;
  assign twiddle4_1_50_imag = T19170 + T19165;
  assign T19165 = {T19168, T19166};
  assign T19166 = $signed(T19167) / $signed(22'h100000);
  assign T19167 = $signed(29'h9c76dd8) * $signed(16'hffff);
  assign T19168 = T19169 ? 2'h3 : 2'h0;
  assign T19169 = T19166[6'h2c:6'h2c];
  assign T19170 = $signed(T19171) / $signed(22'h100000);
  assign T19171 = $signed(31'h3f3f9cab) * $signed(16'h0);
  assign twiddle4_1_51_imag = T19177 + T19172;
  assign T19172 = {T19175, T19173};
  assign T19173 = $signed(T19174) / $signed(22'h100000);
  assign T19174 = $signed(29'h9f917ab) * $signed(16'hffff);
  assign T19175 = T19176 ? 2'h3 : 2'h0;
  assign T19176 = T19173[6'h2c:6'h2c];
  assign T19177 = $signed(T19178) / $signed(22'h100000);
  assign T19178 = $signed(31'h3f37daf9) * $signed(16'h0);
  assign T19179 = T18725[1'h0:1'h0];
  assign T19180 = T18725[1'h1:1'h1];
  assign T19181 = T19214 ? T19198 : T19182;
  assign T19182 = T19197 ? twiddle4_1_53_imag : twiddle4_1_52_imag;
  assign twiddle4_1_52_imag = T19188 + T19183;
  assign T19183 = {T19186, T19184};
  assign T19184 = $signed(T19185) / $signed(22'h100000);
  assign T19185 = $signed(29'ha2abb58) * $signed(16'hffff);
  assign T19186 = T19187 ? 2'h3 : 2'h0;
  assign T19187 = T19184[6'h2c:6'h2c];
  assign T19188 = $signed(T19189) / $signed(22'h100000);
  assign T19189 = $signed(31'h3f2ff249) * $signed(16'h0);
  assign twiddle4_1_53_imag = T19195 + T19190;
  assign T19190 = {T19193, T19191};
  assign T19191 = $signed(T19192) / $signed(22'h100000);
  assign T19192 = $signed(29'ha5c58bf) * $signed(16'hffff);
  assign T19193 = T19194 ? 2'h3 : 2'h0;
  assign T19194 = T19191[6'h2c:6'h2c];
  assign T19195 = $signed(T19196) / $signed(22'h100000);
  assign T19196 = $signed(31'h3f27e29f) * $signed(16'h0);
  assign T19197 = T18725[1'h0:1'h0];
  assign T19198 = T19213 ? twiddle4_1_55_imag : twiddle4_1_54_imag;
  assign twiddle4_1_54_imag = T19204 + T19199;
  assign T19199 = {T19202, T19200};
  assign T19200 = $signed(T19201) / $signed(22'h100000);
  assign T19201 = $signed(29'ha8defc2) * $signed(16'hffff);
  assign T19202 = T19203 ? 2'h3 : 2'h0;
  assign T19203 = T19200[6'h2c:6'h2c];
  assign T19204 = $signed(T19205) / $signed(22'h100000);
  assign T19205 = $signed(31'h3f1fabff) * $signed(16'h0);
  assign twiddle4_1_55_imag = T19211 + T19206;
  assign T19206 = {T19209, T19207};
  assign T19207 = $signed(T19208) / $signed(22'h100000);
  assign T19208 = $signed(29'habf8043) * $signed(16'hffff);
  assign T19209 = T19210 ? 2'h3 : 2'h0;
  assign T19210 = T19207[6'h2c:6'h2c];
  assign T19211 = $signed(T19212) / $signed(22'h100000);
  assign T19212 = $signed(31'h3f174e6f) * $signed(16'h0);
  assign T19213 = T18725[1'h0:1'h0];
  assign T19214 = T18725[1'h1:1'h1];
  assign T19215 = T18725[2'h2:2'h2];
  assign T19216 = T19285 ? T19251 : T19217;
  assign T19217 = T19250 ? T19234 : T19218;
  assign T19218 = T19233 ? twiddle4_1_57_imag : twiddle4_1_56_imag;
  assign twiddle4_1_56_imag = T19224 + T19219;
  assign T19219 = {T19222, T19220};
  assign T19220 = $signed(T19221) / $signed(22'h100000);
  assign T19221 = $signed(29'haf10a22) * $signed(16'hffff);
  assign T19222 = T19223 ? 2'h3 : 2'h0;
  assign T19223 = T19220[6'h2c:6'h2c];
  assign T19224 = $signed(T19225) / $signed(22'h100000);
  assign T19225 = $signed(31'h3f0ec9f4) * $signed(16'h0);
  assign twiddle4_1_57_imag = T19231 + T19226;
  assign T19226 = {T19229, T19227};
  assign T19227 = $signed(T19228) / $signed(22'h100000);
  assign T19228 = $signed(29'hb228d41) * $signed(16'hffff);
  assign T19229 = T19230 ? 2'h3 : 2'h0;
  assign T19230 = T19227[6'h2c:6'h2c];
  assign T19231 = $signed(T19232) / $signed(22'h100000);
  assign T19232 = $signed(31'h3f061e94) * $signed(16'h0);
  assign T19233 = T18725[1'h0:1'h0];
  assign T19234 = T19249 ? twiddle4_1_59_imag : twiddle4_1_58_imag;
  assign twiddle4_1_58_imag = T19240 + T19235;
  assign T19235 = {T19238, T19236};
  assign T19236 = $signed(T19237) / $signed(22'h100000);
  assign T19237 = $signed(29'hb540982) * $signed(16'hffff);
  assign T19238 = T19239 ? 2'h3 : 2'h0;
  assign T19239 = T19236[6'h2c:6'h2c];
  assign T19240 = $signed(T19241) / $signed(22'h100000);
  assign T19241 = $signed(31'h3efd4c53) * $signed(16'h0);
  assign twiddle4_1_59_imag = T19247 + T19242;
  assign T19242 = {T19245, T19243};
  assign T19243 = $signed(T19244) / $signed(22'h100000);
  assign T19244 = $signed(29'hb857ec6) * $signed(16'hffff);
  assign T19245 = T19246 ? 2'h3 : 2'h0;
  assign T19246 = T19243[6'h2c:6'h2c];
  assign T19247 = $signed(T19248) / $signed(22'h100000);
  assign T19248 = $signed(31'h3ef45338) * $signed(16'h0);
  assign T19249 = T18725[1'h0:1'h0];
  assign T19250 = T18725[1'h1:1'h1];
  assign T19251 = T19284 ? T19268 : T19252;
  assign T19252 = T19267 ? twiddle4_1_61_imag : twiddle4_1_60_imag;
  assign twiddle4_1_60_imag = T19258 + T19253;
  assign T19253 = {T19256, T19254};
  assign T19254 = $signed(T19255) / $signed(22'h100000);
  assign T19255 = $signed(29'hbb6ecef) * $signed(16'hffff);
  assign T19256 = T19257 ? 2'h3 : 2'h0;
  assign T19257 = T19254[6'h2c:6'h2c];
  assign T19258 = $signed(T19259) / $signed(22'h100000);
  assign T19259 = $signed(31'h3eeb3347) * $signed(16'h0);
  assign twiddle4_1_61_imag = T19265 + T19260;
  assign T19260 = {T19263, T19261};
  assign T19261 = $signed(T19262) / $signed(22'h100000);
  assign T19262 = $signed(29'hbe853dd) * $signed(16'hffff);
  assign T19263 = T19264 ? 2'h3 : 2'h0;
  assign T19264 = T19261[6'h2c:6'h2c];
  assign T19265 = $signed(T19266) / $signed(22'h100000);
  assign T19266 = $signed(31'h3ee1ec86) * $signed(16'h0);
  assign T19267 = T18725[1'h0:1'h0];
  assign T19268 = T19283 ? twiddle4_1_63_imag : twiddle4_1_62_imag;
  assign twiddle4_1_62_imag = T19274 + T19269;
  assign T19269 = {T19272, T19270};
  assign T19270 = $signed(T19271) / $signed(22'h100000);
  assign T19271 = $signed(29'hc19b374) * $signed(16'hffff);
  assign T19272 = T19273 ? 2'h3 : 2'h0;
  assign T19273 = T19270[6'h2c:6'h2c];
  assign T19274 = $signed(T19275) / $signed(22'h100000);
  assign T19275 = $signed(31'h3ed87efb) * $signed(16'h0);
  assign twiddle4_1_63_imag = T19281 + T19276;
  assign T19276 = {T19279, T19277};
  assign T19277 = $signed(T19278) / $signed(22'h100000);
  assign T19278 = $signed(29'hc4b0b93) * $signed(16'hffff);
  assign T19279 = T19280 ? 2'h3 : 2'h0;
  assign T19280 = T19277[6'h2c:6'h2c];
  assign T19281 = $signed(T19282) / $signed(22'h100000);
  assign T19282 = $signed(31'h3eceeaad) * $signed(16'h0);
  assign T19283 = T18725[1'h0:1'h0];
  assign T19284 = T18725[1'h1:1'h1];
  assign T19285 = T18725[2'h2:2'h2];
  assign T19286 = T18725[2'h3:2'h3];
  assign T19287 = T18725[3'h4:3'h4];
  assign T19288 = T19002[6'h2e:6'h2e];
  assign T19289 = T18725[3'h5:3'h5];
  assign T19290 = {T19820, T19291};
  assign T19291 = T19819 ? T19565 : T19292;
  assign T19292 = T19564 ? T19435 : T19293;
  assign T19293 = T19434 ? T19364 : T19294;
  assign T19294 = T19363 ? T19329 : T19295;
  assign T19295 = T19328 ? T19312 : T19296;
  assign T19296 = T19311 ? twiddle4_1_65_imag : twiddle4_1_64_imag;
  assign twiddle4_1_64_imag = T19302 + T19297;
  assign T19297 = {T19300, T19298};
  assign T19298 = $signed(T19299) / $signed(22'h100000);
  assign T19299 = $signed(29'hc7c5c1e) * $signed(16'hffff);
  assign T19300 = T19301 ? 2'h3 : 2'h0;
  assign T19301 = T19298[6'h2c:6'h2c];
  assign T19302 = $signed(T19303) / $signed(22'h100000);
  assign T19303 = $signed(31'h3ec52f9f) * $signed(16'h0);
  assign twiddle4_1_65_imag = T19309 + T19304;
  assign T19304 = {T19307, T19305};
  assign T19305 = $signed(T19306) / $signed(22'h100000);
  assign T19306 = $signed(29'hcada4f4) * $signed(16'hffff);
  assign T19307 = T19308 ? 2'h3 : 2'h0;
  assign T19308 = T19305[6'h2c:6'h2c];
  assign T19309 = $signed(T19310) / $signed(22'h100000);
  assign T19310 = $signed(31'h3ebb4dda) * $signed(16'h0);
  assign T19311 = T18725[1'h0:1'h0];
  assign T19312 = T19327 ? twiddle4_1_67_imag : twiddle4_1_66_imag;
  assign twiddle4_1_66_imag = T19318 + T19313;
  assign T19313 = {T19316, T19314};
  assign T19314 = $signed(T19315) / $signed(22'h100000);
  assign T19315 = $signed(29'hcdee5f9) * $signed(16'hffff);
  assign T19316 = T19317 ? 2'h3 : 2'h0;
  assign T19317 = T19314[6'h2c:6'h2c];
  assign T19318 = $signed(T19319) / $signed(22'h100000);
  assign T19319 = $signed(31'h3eb14562) * $signed(16'h0);
  assign twiddle4_1_67_imag = T19325 + T19320;
  assign T19320 = {T19323, T19321};
  assign T19321 = $signed(T19322) / $signed(22'h100000);
  assign T19322 = $signed(29'hd101f0d) * $signed(16'hffff);
  assign T19323 = T19324 ? 2'h3 : 2'h0;
  assign T19324 = T19321[6'h2c:6'h2c];
  assign T19325 = $signed(T19326) / $signed(22'h100000);
  assign T19326 = $signed(31'h3ea7163f) * $signed(16'h0);
  assign T19327 = T18725[1'h0:1'h0];
  assign T19328 = T18725[1'h1:1'h1];
  assign T19329 = T19362 ? T19346 : T19330;
  assign T19330 = T19345 ? twiddle4_1_69_imag : twiddle4_1_68_imag;
  assign twiddle4_1_68_imag = T19336 + T19331;
  assign T19331 = {T19334, T19332};
  assign T19332 = $signed(T19333) / $signed(22'h100000);
  assign T19333 = $signed(29'hd415012) * $signed(16'hffff);
  assign T19334 = T19335 ? 2'h3 : 2'h0;
  assign T19335 = T19332[6'h2c:6'h2c];
  assign T19336 = $signed(T19337) / $signed(22'h100000);
  assign T19337 = $signed(31'h3e9cc076) * $signed(16'h0);
  assign twiddle4_1_69_imag = T19343 + T19338;
  assign T19338 = {T19341, T19339};
  assign T19339 = $signed(T19340) / $signed(22'h100000);
  assign T19340 = $signed(29'hd7278ea) * $signed(16'hffff);
  assign T19341 = T19342 ? 2'h3 : 2'h0;
  assign T19342 = T19339[6'h2c:6'h2c];
  assign T19343 = $signed(T19344) / $signed(22'h100000);
  assign T19344 = $signed(31'h3e92440d) * $signed(16'h0);
  assign T19345 = T18725[1'h0:1'h0];
  assign T19346 = T19361 ? twiddle4_1_71_imag : twiddle4_1_70_imag;
  assign twiddle4_1_70_imag = T19352 + T19347;
  assign T19347 = {T19350, T19348};
  assign T19348 = $signed(T19349) / $signed(22'h100000);
  assign T19349 = $signed(29'hda39977) * $signed(16'hffff);
  assign T19350 = T19351 ? 2'h3 : 2'h0;
  assign T19351 = T19348[6'h2c:6'h2c];
  assign T19352 = $signed(T19353) / $signed(22'h100000);
  assign T19353 = $signed(31'h3e87a10b) * $signed(16'h0);
  assign twiddle4_1_71_imag = T19359 + T19354;
  assign T19354 = {T19357, T19355};
  assign T19355 = $signed(T19356) / $signed(22'h100000);
  assign T19356 = $signed(29'hdd4b19a) * $signed(16'hffff);
  assign T19357 = T19358 ? 2'h3 : 2'h0;
  assign T19358 = T19355[6'h2c:6'h2c];
  assign T19359 = $signed(T19360) / $signed(22'h100000);
  assign T19360 = $signed(31'h3e7cd778) * $signed(16'h0);
  assign T19361 = T18725[1'h0:1'h0];
  assign T19362 = T18725[1'h1:1'h1];
  assign T19363 = T18725[2'h2:2'h2];
  assign T19364 = T19433 ? T19399 : T19365;
  assign T19365 = T19398 ? T19382 : T19366;
  assign T19366 = T19381 ? twiddle4_1_73_imag : twiddle4_1_72_imag;
  assign twiddle4_1_72_imag = T19372 + T19367;
  assign T19367 = {T19370, T19368};
  assign T19368 = $signed(T19369) / $signed(22'h100000);
  assign T19369 = $signed(29'he05c135) * $signed(16'hffff);
  assign T19370 = T19371 ? 2'h3 : 2'h0;
  assign T19371 = T19368[6'h2c:6'h2c];
  assign T19372 = $signed(T19373) / $signed(22'h100000);
  assign T19373 = $signed(31'h3e71e758) * $signed(16'h0);
  assign twiddle4_1_73_imag = T19379 + T19374;
  assign T19374 = {T19377, T19375};
  assign T19375 = $signed(T19376) / $signed(22'h100000);
  assign T19376 = $signed(29'he36c829) * $signed(16'hffff);
  assign T19377 = T19378 ? 2'h3 : 2'h0;
  assign T19378 = T19375[6'h2c:6'h2c];
  assign T19379 = $signed(T19380) / $signed(22'h100000);
  assign T19380 = $signed(31'h3e66d0b4) * $signed(16'h0);
  assign T19381 = T18725[1'h0:1'h0];
  assign T19382 = T19397 ? twiddle4_1_75_imag : twiddle4_1_74_imag;
  assign twiddle4_1_74_imag = T19388 + T19383;
  assign T19383 = {T19386, T19384};
  assign T19384 = $signed(T19385) / $signed(22'h100000);
  assign T19385 = $signed(29'he67c659) * $signed(16'hffff);
  assign T19386 = T19387 ? 2'h3 : 2'h0;
  assign T19387 = T19384[6'h2c:6'h2c];
  assign T19388 = $signed(T19389) / $signed(22'h100000);
  assign T19389 = $signed(31'h3e5b9392) * $signed(16'h0);
  assign twiddle4_1_75_imag = T19395 + T19390;
  assign T19390 = {T19393, T19391};
  assign T19391 = $signed(T19392) / $signed(22'h100000);
  assign T19392 = $signed(29'he98bba6) * $signed(16'hffff);
  assign T19393 = T19394 ? 2'h3 : 2'h0;
  assign T19394 = T19391[6'h2c:6'h2c];
  assign T19395 = $signed(T19396) / $signed(22'h100000);
  assign T19396 = $signed(31'h3e502ff8) * $signed(16'h0);
  assign T19397 = T18725[1'h0:1'h0];
  assign T19398 = T18725[1'h1:1'h1];
  assign T19399 = T19432 ? T19416 : T19400;
  assign T19400 = T19415 ? twiddle4_1_77_imag : twiddle4_1_76_imag;
  assign twiddle4_1_76_imag = T19406 + T19401;
  assign T19401 = {T19404, T19402};
  assign T19402 = $signed(T19403) / $signed(22'h100000);
  assign T19403 = $signed(29'hec9a7f2) * $signed(16'hffff);
  assign T19404 = T19405 ? 2'h3 : 2'h0;
  assign T19405 = T19402[6'h2c:6'h2c];
  assign T19406 = $signed(T19407) / $signed(22'h100000);
  assign T19407 = $signed(31'h3e44a5ee) * $signed(16'h0);
  assign twiddle4_1_77_imag = T19413 + T19408;
  assign T19408 = {T19411, T19409};
  assign T19409 = $signed(T19410) / $signed(22'h100000);
  assign T19410 = $signed(29'hefa8b1f) * $signed(16'hffff);
  assign T19411 = T19412 ? 2'h3 : 2'h0;
  assign T19412 = T19409[6'h2c:6'h2c];
  assign T19413 = $signed(T19414) / $signed(22'h100000);
  assign T19414 = $signed(31'h3e38f57c) * $signed(16'h0);
  assign T19415 = T18725[1'h0:1'h0];
  assign T19416 = T19431 ? twiddle4_1_79_imag : twiddle4_1_78_imag;
  assign twiddle4_1_78_imag = T19422 + T19417;
  assign T19417 = {T19420, T19418};
  assign T19418 = $signed(T19419) / $signed(22'h100000);
  assign T19419 = $signed(29'hf2b650f) * $signed(16'hffff);
  assign T19420 = T19421 ? 2'h3 : 2'h0;
  assign T19421 = T19418[6'h2c:6'h2c];
  assign T19422 = $signed(T19423) / $signed(22'h100000);
  assign T19423 = $signed(31'h3e2d1ea7) * $signed(16'h0);
  assign twiddle4_1_79_imag = T19429 + T19424;
  assign T19424 = {T19427, T19425};
  assign T19425 = $signed(T19426) / $signed(22'h100000);
  assign T19426 = $signed(29'hf5c35a3) * $signed(16'hffff);
  assign T19427 = T19428 ? 2'h3 : 2'h0;
  assign T19428 = T19425[6'h2c:6'h2c];
  assign T19429 = $signed(T19430) / $signed(22'h100000);
  assign T19430 = $signed(31'h3e212179) * $signed(16'h0);
  assign T19431 = T18725[1'h0:1'h0];
  assign T19432 = T18725[1'h1:1'h1];
  assign T19433 = T18725[2'h2:2'h2];
  assign T19434 = T18725[2'h3:2'h3];
  assign T19435 = T19563 ? T19501 : T19436;
  assign T19436 = T19500 ? T19470 : T19437;
  assign T19437 = T19469 ? T19454 : T19438;
  assign T19438 = T19453 ? twiddle4_1_81_imag : twiddle4_1_80_imag;
  assign twiddle4_1_80_imag = T19444 + T19439;
  assign T19439 = {T19442, T19440};
  assign T19440 = $signed(T19441) / $signed(22'h100000);
  assign T19441 = $signed(29'hf8cfcbd) * $signed(16'hffff);
  assign T19442 = T19443 ? 2'h3 : 2'h0;
  assign T19443 = T19440[6'h2c:6'h2c];
  assign T19444 = $signed(T19445) / $signed(22'h100000);
  assign T19445 = $signed(31'h3e14fdf7) * $signed(16'h0);
  assign twiddle4_1_81_imag = T19451 + T19446;
  assign T19446 = {T19449, T19447};
  assign T19447 = $signed(T19448) / $signed(22'h100000);
  assign T19448 = $signed(29'hfbdba40) * $signed(16'hffff);
  assign T19449 = T19450 ? 2'h3 : 2'h0;
  assign T19450 = T19447[6'h2c:6'h2c];
  assign T19451 = $signed(T19452) / $signed(22'h100000);
  assign T19452 = $signed(31'h3e08b429) * $signed(16'h0);
  assign T19453 = T18725[1'h0:1'h0];
  assign T19454 = T19468 ? twiddle4_1_83_imag : twiddle4_1_82_imag;
  assign twiddle4_1_82_imag = T19460 + T19455;
  assign T19455 = {T19458, T19456};
  assign T19456 = $signed(T19457) / $signed(22'h100000);
  assign T19457 = $signed(29'hfee6e0d) * $signed(16'hffff);
  assign T19458 = T19459 ? 2'h3 : 2'h0;
  assign T19459 = T19456[6'h2c:6'h2c];
  assign T19460 = $signed(T19461) / $signed(22'h100000);
  assign T19461 = $signed(31'h3dfc4418) * $signed(16'h0);
  assign twiddle4_1_83_imag = T19466 + T19462;
  assign T19462 = {T19465, T19463};
  assign T19463 = $signed(T19464) / $signed(22'h100000);
  assign T19464 = $signed(30'h101f1806) * $signed(16'hffff);
  assign T19465 = T19463[6'h2d:6'h2d];
  assign T19466 = $signed(T19467) / $signed(22'h100000);
  assign T19467 = $signed(31'h3defadca) * $signed(16'h0);
  assign T19468 = T18725[1'h0:1'h0];
  assign T19469 = T18725[1'h1:1'h1];
  assign T19470 = T19499 ? T19485 : T19471;
  assign T19471 = T19484 ? twiddle4_1_85_imag : twiddle4_1_84_imag;
  assign twiddle4_1_84_imag = T19476 + T19472;
  assign T19472 = {T19475, T19473};
  assign T19473 = $signed(T19474) / $signed(22'h100000);
  assign T19474 = $signed(30'h104fb80e) * $signed(16'hffff);
  assign T19475 = T19473[6'h2d:6'h2d];
  assign T19476 = $signed(T19477) / $signed(22'h100000);
  assign T19477 = $signed(31'h3de2f147) * $signed(16'h0);
  assign twiddle4_1_85_imag = T19482 + T19478;
  assign T19478 = {T19481, T19479};
  assign T19479 = $signed(T19480) / $signed(22'h100000);
  assign T19480 = $signed(30'h10804e05) * $signed(16'hffff);
  assign T19481 = T19479[6'h2d:6'h2d];
  assign T19482 = $signed(T19483) / $signed(22'h100000);
  assign T19483 = $signed(31'h3dd60e98) * $signed(16'h0);
  assign T19484 = T18725[1'h0:1'h0];
  assign T19485 = T19498 ? twiddle4_1_87_imag : twiddle4_1_86_imag;
  assign twiddle4_1_86_imag = T19490 + T19486;
  assign T19486 = {T19489, T19487};
  assign T19487 = $signed(T19488) / $signed(22'h100000);
  assign T19488 = $signed(30'h10b0d9cf) * $signed(16'hffff);
  assign T19489 = T19487[6'h2d:6'h2d];
  assign T19490 = $signed(T19491) / $signed(22'h100000);
  assign T19491 = $signed(31'h3dc905c4) * $signed(16'h0);
  assign twiddle4_1_87_imag = T19496 + T19492;
  assign T19492 = {T19495, T19493};
  assign T19493 = $signed(T19494) / $signed(22'h100000);
  assign T19494 = $signed(30'h10e15b4e) * $signed(16'hffff);
  assign T19495 = T19493[6'h2d:6'h2d];
  assign T19496 = $signed(T19497) / $signed(22'h100000);
  assign T19497 = $signed(31'h3dbbd6d4) * $signed(16'h0);
  assign T19498 = T18725[1'h0:1'h0];
  assign T19499 = T18725[1'h1:1'h1];
  assign T19500 = T18725[2'h2:2'h2];
  assign T19501 = T19562 ? T19532 : T19502;
  assign T19502 = T19531 ? T19517 : T19503;
  assign T19503 = T19516 ? twiddle4_1_89_imag : twiddle4_1_88_imag;
  assign twiddle4_1_88_imag = T19508 + T19504;
  assign T19504 = {T19507, T19505};
  assign T19505 = $signed(T19506) / $signed(22'h100000);
  assign T19506 = $signed(30'h1111d262) * $signed(16'hffff);
  assign T19507 = T19505[6'h2d:6'h2d];
  assign T19508 = $signed(T19509) / $signed(22'h100000);
  assign T19509 = $signed(31'h3dae81ce) * $signed(16'h0);
  assign twiddle4_1_89_imag = T19514 + T19510;
  assign T19510 = {T19513, T19511};
  assign T19511 = $signed(T19512) / $signed(22'h100000);
  assign T19512 = $signed(30'h11423eef) * $signed(16'hffff);
  assign T19513 = T19511[6'h2d:6'h2d];
  assign T19514 = $signed(T19515) / $signed(22'h100000);
  assign T19515 = $signed(31'h3da106bd) * $signed(16'h0);
  assign T19516 = T18725[1'h0:1'h0];
  assign T19517 = T19530 ? twiddle4_1_91_imag : twiddle4_1_90_imag;
  assign twiddle4_1_90_imag = T19522 + T19518;
  assign T19518 = {T19521, T19519};
  assign T19519 = $signed(T19520) / $signed(22'h100000);
  assign T19520 = $signed(30'h1172a0d7) * $signed(16'hffff);
  assign T19521 = T19519[6'h2d:6'h2d];
  assign T19522 = $signed(T19523) / $signed(22'h100000);
  assign T19523 = $signed(31'h3d9365a7) * $signed(16'h0);
  assign twiddle4_1_91_imag = T19528 + T19524;
  assign T19524 = {T19527, T19525};
  assign T19525 = $signed(T19526) / $signed(22'h100000);
  assign T19526 = $signed(30'h11a2f7fb) * $signed(16'hffff);
  assign T19527 = T19525[6'h2d:6'h2d];
  assign T19528 = $signed(T19529) / $signed(22'h100000);
  assign T19529 = $signed(31'h3d859e96) * $signed(16'h0);
  assign T19530 = T18725[1'h0:1'h0];
  assign T19531 = T18725[1'h1:1'h1];
  assign T19532 = T19561 ? T19547 : T19533;
  assign T19533 = T19546 ? twiddle4_1_93_imag : twiddle4_1_92_imag;
  assign twiddle4_1_92_imag = T19538 + T19534;
  assign T19534 = {T19537, T19535};
  assign T19535 = $signed(T19536) / $signed(22'h100000);
  assign T19536 = $signed(30'h11d3443f) * $signed(16'hffff);
  assign T19537 = T19535[6'h2d:6'h2d];
  assign T19538 = $signed(T19539) / $signed(22'h100000);
  assign T19539 = $signed(31'h3d77b191) * $signed(16'h0);
  assign twiddle4_1_93_imag = T19544 + T19540;
  assign T19540 = {T19543, T19541};
  assign T19541 = $signed(T19542) / $signed(22'h100000);
  assign T19542 = $signed(30'h12038583) * $signed(16'hffff);
  assign T19543 = T19541[6'h2d:6'h2d];
  assign T19544 = $signed(T19545) / $signed(22'h100000);
  assign T19545 = $signed(31'h3d699ea2) * $signed(16'h0);
  assign T19546 = T18725[1'h0:1'h0];
  assign T19547 = T19560 ? twiddle4_1_95_imag : twiddle4_1_94_imag;
  assign twiddle4_1_94_imag = T19552 + T19548;
  assign T19548 = {T19551, T19549};
  assign T19549 = $signed(T19550) / $signed(22'h100000);
  assign T19550 = $signed(30'h1233bbab) * $signed(16'hffff);
  assign T19551 = T19549[6'h2d:6'h2d];
  assign T19552 = $signed(T19553) / $signed(22'h100000);
  assign T19553 = $signed(31'h3d5b65d1) * $signed(16'h0);
  assign twiddle4_1_95_imag = T19558 + T19554;
  assign T19554 = {T19557, T19555};
  assign T19555 = $signed(T19556) / $signed(22'h100000);
  assign T19556 = $signed(30'h1263e699) * $signed(16'hffff);
  assign T19557 = T19555[6'h2d:6'h2d];
  assign T19558 = $signed(T19559) / $signed(22'h100000);
  assign T19559 = $signed(31'h3d4d0727) * $signed(16'h0);
  assign T19560 = T18725[1'h0:1'h0];
  assign T19561 = T18725[1'h1:1'h1];
  assign T19562 = T18725[2'h2:2'h2];
  assign T19563 = T18725[2'h3:2'h3];
  assign T19564 = T18725[3'h4:3'h4];
  assign T19565 = T19818 ? T19692 : T19566;
  assign T19566 = T19691 ? T19629 : T19567;
  assign T19567 = T19628 ? T19598 : T19568;
  assign T19568 = T19597 ? T19583 : T19569;
  assign T19569 = T19582 ? twiddle4_1_97_imag : twiddle4_1_96_imag;
  assign twiddle4_1_96_imag = T19574 + T19570;
  assign T19570 = {T19573, T19571};
  assign T19571 = $signed(T19572) / $signed(22'h100000);
  assign T19572 = $signed(30'h1294062e) * $signed(16'hffff);
  assign T19573 = T19571[6'h2d:6'h2d];
  assign T19574 = $signed(T19575) / $signed(22'h100000);
  assign T19575 = $signed(31'h3d3e82ad) * $signed(16'h0);
  assign twiddle4_1_97_imag = T19580 + T19576;
  assign T19576 = {T19579, T19577};
  assign T19577 = $signed(T19578) / $signed(22'h100000);
  assign T19578 = $signed(30'h12c41a4e) * $signed(16'hffff);
  assign T19579 = T19577[6'h2d:6'h2d];
  assign T19580 = $signed(T19581) / $signed(22'h100000);
  assign T19581 = $signed(31'h3d2fd86c) * $signed(16'h0);
  assign T19582 = T18725[1'h0:1'h0];
  assign T19583 = T19596 ? twiddle4_1_99_imag : twiddle4_1_98_imag;
  assign twiddle4_1_98_imag = T19588 + T19584;
  assign T19584 = {T19587, T19585};
  assign T19585 = $signed(T19586) / $signed(22'h100000);
  assign T19586 = $signed(30'h12f422da) * $signed(16'hffff);
  assign T19587 = T19585[6'h2d:6'h2d];
  assign T19588 = $signed(T19589) / $signed(22'h100000);
  assign T19589 = $signed(31'h3d21086c) * $signed(16'h0);
  assign twiddle4_1_99_imag = T19594 + T19590;
  assign T19590 = {T19593, T19591};
  assign T19591 = $signed(T19592) / $signed(22'h100000);
  assign T19592 = $signed(30'h13241fb6) * $signed(16'hffff);
  assign T19593 = T19591[6'h2d:6'h2d];
  assign T19594 = $signed(T19595) / $signed(22'h100000);
  assign T19595 = $signed(31'h3d1212b7) * $signed(16'h0);
  assign T19596 = T18725[1'h0:1'h0];
  assign T19597 = T18725[1'h1:1'h1];
  assign T19598 = T19627 ? T19613 : T19599;
  assign T19599 = T19612 ? twiddle4_1_101_imag : twiddle4_1_100_imag;
  assign twiddle4_1_100_imag = T19604 + T19600;
  assign T19600 = {T19603, T19601};
  assign T19601 = $signed(T19602) / $signed(22'h100000);
  assign T19602 = $signed(30'h135410c2) * $signed(16'hffff);
  assign T19603 = T19601[6'h2d:6'h2d];
  assign T19604 = $signed(T19605) / $signed(22'h100000);
  assign T19605 = $signed(31'h3d02f756) * $signed(16'h0);
  assign twiddle4_1_101_imag = T19610 + T19606;
  assign T19606 = {T19609, T19607};
  assign T19607 = $signed(T19608) / $signed(22'h100000);
  assign T19608 = $signed(30'h1383f5e3) * $signed(16'hffff);
  assign T19609 = T19607[6'h2d:6'h2d];
  assign T19610 = $signed(T19611) / $signed(22'h100000);
  assign T19611 = $signed(31'h3cf3b653) * $signed(16'h0);
  assign T19612 = T18725[1'h0:1'h0];
  assign T19613 = T19626 ? twiddle4_1_103_imag : twiddle4_1_102_imag;
  assign twiddle4_1_102_imag = T19618 + T19614;
  assign T19614 = {T19617, T19615};
  assign T19615 = $signed(T19616) / $signed(22'h100000);
  assign T19616 = $signed(30'h13b3cefa) * $signed(16'hffff);
  assign T19617 = T19615[6'h2d:6'h2d];
  assign T19618 = $signed(T19619) / $signed(22'h100000);
  assign T19619 = $signed(31'h3ce44fb6) * $signed(16'h0);
  assign twiddle4_1_103_imag = T19624 + T19620;
  assign T19620 = {T19623, T19621};
  assign T19621 = $signed(T19622) / $signed(22'h100000);
  assign T19622 = $signed(30'h13e39be9) * $signed(16'hffff);
  assign T19623 = T19621[6'h2d:6'h2d];
  assign T19624 = $signed(T19625) / $signed(22'h100000);
  assign T19625 = $signed(31'h3cd4c38a) * $signed(16'h0);
  assign T19626 = T18725[1'h0:1'h0];
  assign T19627 = T18725[1'h1:1'h1];
  assign T19628 = T18725[2'h2:2'h2];
  assign T19629 = T19690 ? T19660 : T19630;
  assign T19630 = T19659 ? T19645 : T19631;
  assign T19631 = T19644 ? twiddle4_1_105_imag : twiddle4_1_104_imag;
  assign twiddle4_1_104_imag = T19636 + T19632;
  assign T19632 = {T19635, T19633};
  assign T19633 = $signed(T19634) / $signed(22'h100000);
  assign T19634 = $signed(30'h14135c94) * $signed(16'hffff);
  assign T19635 = T19633[6'h2d:6'h2d];
  assign T19636 = $signed(T19637) / $signed(22'h100000);
  assign T19637 = $signed(31'h3cc511d8) * $signed(16'h0);
  assign twiddle4_1_105_imag = T19642 + T19638;
  assign T19638 = {T19641, T19639};
  assign T19639 = $signed(T19640) / $signed(22'h100000);
  assign T19640 = $signed(30'h144310dc) * $signed(16'hffff);
  assign T19641 = T19639[6'h2d:6'h2d];
  assign T19642 = $signed(T19643) / $signed(22'h100000);
  assign T19643 = $signed(31'h3cb53aaa) * $signed(16'h0);
  assign T19644 = T18725[1'h0:1'h0];
  assign T19645 = T19658 ? twiddle4_1_107_imag : twiddle4_1_106_imag;
  assign twiddle4_1_106_imag = T19650 + T19646;
  assign T19646 = {T19649, T19647};
  assign T19647 = $signed(T19648) / $signed(22'h100000);
  assign T19648 = $signed(30'h1472b8a5) * $signed(16'hffff);
  assign T19649 = T19647[6'h2d:6'h2d];
  assign T19650 = $signed(T19651) / $signed(22'h100000);
  assign T19651 = $signed(31'h3ca53e08) * $signed(16'h0);
  assign twiddle4_1_107_imag = T19656 + T19652;
  assign T19652 = {T19655, T19653};
  assign T19653 = $signed(T19654) / $signed(22'h100000);
  assign T19654 = $signed(30'h14a253d1) * $signed(16'hffff);
  assign T19655 = T19653[6'h2d:6'h2d];
  assign T19656 = $signed(T19657) / $signed(22'h100000);
  assign T19657 = $signed(31'h3c951bff) * $signed(16'h0);
  assign T19658 = T18725[1'h0:1'h0];
  assign T19659 = T18725[1'h1:1'h1];
  assign T19660 = T19689 ? T19675 : T19661;
  assign T19661 = T19674 ? twiddle4_1_109_imag : twiddle4_1_108_imag;
  assign twiddle4_1_108_imag = T19666 + T19662;
  assign T19662 = {T19665, T19663};
  assign T19663 = $signed(T19664) / $signed(22'h100000);
  assign T19664 = $signed(30'h14d1e242) * $signed(16'hffff);
  assign T19665 = T19663[6'h2d:6'h2d];
  assign T19666 = $signed(T19667) / $signed(22'h100000);
  assign T19667 = $signed(31'h3c84d496) * $signed(16'h0);
  assign twiddle4_1_109_imag = T19672 + T19668;
  assign T19668 = {T19671, T19669};
  assign T19669 = $signed(T19670) / $signed(22'h100000);
  assign T19670 = $signed(30'h150163dc) * $signed(16'hffff);
  assign T19671 = T19669[6'h2d:6'h2d];
  assign T19672 = $signed(T19673) / $signed(22'h100000);
  assign T19673 = $signed(31'h3c7467d8) * $signed(16'h0);
  assign T19674 = T18725[1'h0:1'h0];
  assign T19675 = T19688 ? twiddle4_1_111_imag : twiddle4_1_110_imag;
  assign twiddle4_1_110_imag = T19680 + T19676;
  assign T19676 = {T19679, T19677};
  assign T19677 = $signed(T19678) / $signed(22'h100000);
  assign T19678 = $signed(30'h1530d880) * $signed(16'hffff);
  assign T19679 = T19677[6'h2d:6'h2d];
  assign T19680 = $signed(T19681) / $signed(22'h100000);
  assign T19681 = $signed(31'h3c63d5d0) * $signed(16'h0);
  assign twiddle4_1_111_imag = T19686 + T19682;
  assign T19682 = {T19685, T19683};
  assign T19683 = $signed(T19684) / $signed(22'h100000);
  assign T19684 = $signed(30'h15604012) * $signed(16'hffff);
  assign T19685 = T19683[6'h2d:6'h2d];
  assign T19686 = $signed(T19687) / $signed(22'h100000);
  assign T19687 = $signed(31'h3c531e88) * $signed(16'h0);
  assign T19688 = T18725[1'h0:1'h0];
  assign T19689 = T18725[1'h1:1'h1];
  assign T19690 = T18725[2'h2:2'h2];
  assign T19691 = T18725[2'h3:2'h3];
  assign T19692 = T19817 ? T19755 : T19693;
  assign T19693 = T19754 ? T19724 : T19694;
  assign T19694 = T19723 ? T19709 : T19695;
  assign T19695 = T19708 ? twiddle4_1_113_imag : twiddle4_1_112_imag;
  assign twiddle4_1_112_imag = T19700 + T19696;
  assign T19696 = {T19699, T19697};
  assign T19697 = $signed(T19698) / $signed(22'h100000);
  assign T19698 = $signed(30'h158f9a75) * $signed(16'hffff);
  assign T19699 = T19697[6'h2d:6'h2d];
  assign T19700 = $signed(T19701) / $signed(22'h100000);
  assign T19701 = $signed(31'h3c424209) * $signed(16'h0);
  assign twiddle4_1_113_imag = T19706 + T19702;
  assign T19702 = {T19705, T19703};
  assign T19703 = $signed(T19704) / $signed(22'h100000);
  assign T19704 = $signed(30'h15bee78b) * $signed(16'hffff);
  assign T19705 = T19703[6'h2d:6'h2d];
  assign T19706 = $signed(T19707) / $signed(22'h100000);
  assign T19707 = $signed(31'h3c31405f) * $signed(16'h0);
  assign T19708 = T18725[1'h0:1'h0];
  assign T19709 = T19722 ? twiddle4_1_115_imag : twiddle4_1_114_imag;
  assign twiddle4_1_114_imag = T19714 + T19710;
  assign T19710 = {T19713, T19711};
  assign T19711 = $signed(T19712) / $signed(22'h100000);
  assign T19712 = $signed(30'h15ee2737) * $signed(16'hffff);
  assign T19713 = T19711[6'h2d:6'h2d];
  assign T19714 = $signed(T19715) / $signed(22'h100000);
  assign T19715 = $signed(31'h3c201994) * $signed(16'h0);
  assign twiddle4_1_115_imag = T19720 + T19716;
  assign T19716 = {T19719, T19717};
  assign T19717 = $signed(T19718) / $signed(22'h100000);
  assign T19718 = $signed(30'h161d595c) * $signed(16'hffff);
  assign T19719 = T19717[6'h2d:6'h2d];
  assign T19720 = $signed(T19721) / $signed(22'h100000);
  assign T19721 = $signed(31'h3c0ecdb2) * $signed(16'h0);
  assign T19722 = T18725[1'h0:1'h0];
  assign T19723 = T18725[1'h1:1'h1];
  assign T19724 = T19753 ? T19739 : T19725;
  assign T19725 = T19738 ? twiddle4_1_117_imag : twiddle4_1_116_imag;
  assign twiddle4_1_116_imag = T19730 + T19726;
  assign T19726 = {T19729, T19727};
  assign T19727 = $signed(T19728) / $signed(22'h100000);
  assign T19728 = $signed(30'h164c7ddd) * $signed(16'hffff);
  assign T19729 = T19727[6'h2d:6'h2d];
  assign T19730 = $signed(T19731) / $signed(22'h100000);
  assign T19731 = $signed(31'h3bfd5cc4) * $signed(16'h0);
  assign twiddle4_1_117_imag = T19736 + T19732;
  assign T19732 = {T19735, T19733};
  assign T19733 = $signed(T19734) / $signed(22'h100000);
  assign T19734 = $signed(30'h167b949c) * $signed(16'hffff);
  assign T19735 = T19733[6'h2d:6'h2d];
  assign T19736 = $signed(T19737) / $signed(22'h100000);
  assign T19737 = $signed(31'h3bebc6d5) * $signed(16'h0);
  assign T19738 = T18725[1'h0:1'h0];
  assign T19739 = T19752 ? twiddle4_1_119_imag : twiddle4_1_118_imag;
  assign twiddle4_1_118_imag = T19744 + T19740;
  assign T19740 = {T19743, T19741};
  assign T19741 = $signed(T19742) / $signed(22'h100000);
  assign T19742 = $signed(30'h16aa9d7d) * $signed(16'hffff);
  assign T19743 = T19741[6'h2d:6'h2d];
  assign T19744 = $signed(T19745) / $signed(22'h100000);
  assign T19745 = $signed(31'h3bda0bef) * $signed(16'h0);
  assign twiddle4_1_119_imag = T19750 + T19746;
  assign T19746 = {T19749, T19747};
  assign T19747 = $signed(T19748) / $signed(22'h100000);
  assign T19748 = $signed(30'h16d99863) * $signed(16'hffff);
  assign T19749 = T19747[6'h2d:6'h2d];
  assign T19750 = $signed(T19751) / $signed(22'h100000);
  assign T19751 = $signed(31'h3bc82c1e) * $signed(16'h0);
  assign T19752 = T18725[1'h0:1'h0];
  assign T19753 = T18725[1'h1:1'h1];
  assign T19754 = T18725[2'h2:2'h2];
  assign T19755 = T19816 ? T19786 : T19756;
  assign T19756 = T19785 ? T19771 : T19757;
  assign T19757 = T19770 ? twiddle4_1_121_imag : twiddle4_1_120_imag;
  assign twiddle4_1_120_imag = T19762 + T19758;
  assign T19758 = {T19761, T19759};
  assign T19759 = $signed(T19760) / $signed(22'h100000);
  assign T19760 = $signed(30'h17088530) * $signed(16'hffff);
  assign T19761 = T19759[6'h2d:6'h2d];
  assign T19762 = $signed(T19763) / $signed(22'h100000);
  assign T19763 = $signed(31'h3bb6276d) * $signed(16'h0);
  assign twiddle4_1_121_imag = T19768 + T19764;
  assign T19764 = {T19767, T19765};
  assign T19765 = $signed(T19766) / $signed(22'h100000);
  assign T19766 = $signed(30'h173763c9) * $signed(16'hffff);
  assign T19767 = T19765[6'h2d:6'h2d];
  assign T19768 = $signed(T19769) / $signed(22'h100000);
  assign T19769 = $signed(31'h3ba3fde7) * $signed(16'h0);
  assign T19770 = T18725[1'h0:1'h0];
  assign T19771 = T19784 ? twiddle4_1_123_imag : twiddle4_1_122_imag;
  assign twiddle4_1_122_imag = T19776 + T19772;
  assign T19772 = {T19775, T19773};
  assign T19773 = $signed(T19774) / $signed(22'h100000);
  assign T19774 = $signed(30'h1766340f) * $signed(16'hffff);
  assign T19775 = T19773[6'h2d:6'h2d];
  assign T19776 = $signed(T19777) / $signed(22'h100000);
  assign T19777 = $signed(31'h3b91af96) * $signed(16'h0);
  assign twiddle4_1_123_imag = T19782 + T19778;
  assign T19778 = {T19781, T19779};
  assign T19779 = $signed(T19780) / $signed(22'h100000);
  assign T19780 = $signed(30'h1794f5e6) * $signed(16'hffff);
  assign T19781 = T19779[6'h2d:6'h2d];
  assign T19782 = $signed(T19783) / $signed(22'h100000);
  assign T19783 = $signed(31'h3b7f3c87) * $signed(16'h0);
  assign T19784 = T18725[1'h0:1'h0];
  assign T19785 = T18725[1'h1:1'h1];
  assign T19786 = T19815 ? T19801 : T19787;
  assign T19787 = T19800 ? twiddle4_1_125_imag : twiddle4_1_124_imag;
  assign twiddle4_1_124_imag = T19792 + T19788;
  assign T19788 = {T19791, T19789};
  assign T19789 = $signed(T19790) / $signed(22'h100000);
  assign T19790 = $signed(30'h17c3a931) * $signed(16'hffff);
  assign T19791 = T19789[6'h2d:6'h2d];
  assign T19792 = $signed(T19793) / $signed(22'h100000);
  assign T19793 = $signed(31'h3b6ca4c4) * $signed(16'h0);
  assign twiddle4_1_125_imag = T19798 + T19794;
  assign T19794 = {T19797, T19795};
  assign T19795 = $signed(T19796) / $signed(22'h100000);
  assign T19796 = $signed(30'h17f24dd3) * $signed(16'hffff);
  assign T19797 = T19795[6'h2d:6'h2d];
  assign T19798 = $signed(T19799) / $signed(22'h100000);
  assign T19799 = $signed(31'h3b59e859) * $signed(16'h0);
  assign T19800 = T18725[1'h0:1'h0];
  assign T19801 = T19814 ? twiddle4_1_127_imag : twiddle4_1_126_imag;
  assign twiddle4_1_126_imag = T19806 + T19802;
  assign T19802 = {T19805, T19803};
  assign T19803 = $signed(T19804) / $signed(22'h100000);
  assign T19804 = $signed(30'h1820e3b0) * $signed(16'hffff);
  assign T19805 = T19803[6'h2d:6'h2d];
  assign T19806 = $signed(T19807) / $signed(22'h100000);
  assign T19807 = $signed(31'h3b470752) * $signed(16'h0);
  assign twiddle4_1_127_imag = T19812 + T19808;
  assign T19808 = {T19811, T19809};
  assign T19809 = $signed(T19810) / $signed(22'h100000);
  assign T19810 = $signed(30'h184f6aaa) * $signed(16'hffff);
  assign T19811 = T19809[6'h2d:6'h2d];
  assign T19812 = $signed(T19813) / $signed(22'h100000);
  assign T19813 = $signed(31'h3b3401bb) * $signed(16'h0);
  assign T19814 = T18725[1'h0:1'h0];
  assign T19815 = T18725[1'h1:1'h1];
  assign T19816 = T18725[2'h2:2'h2];
  assign T19817 = T18725[2'h3:2'h3];
  assign T19818 = T18725[3'h4:3'h4];
  assign T19819 = T18725[3'h5:3'h5];
  assign T19820 = T19291[6'h2e:6'h2e];
  assign T19821 = T18725[3'h6:3'h6];
  assign T19822 = {T20675, T19823};
  assign T19823 = T20674 ? T20292 : T19824;
  assign T19824 = T20291 ? T20079 : T19825;
  assign T19825 = T20078 ? T19952 : T19826;
  assign T19826 = T19951 ? T19889 : T19827;
  assign T19827 = T19888 ? T19858 : T19828;
  assign T19828 = T19857 ? T19843 : T19829;
  assign T19829 = T19842 ? twiddle4_1_129_imag : twiddle4_1_128_imag;
  assign twiddle4_1_128_imag = T19834 + T19830;
  assign T19830 = {T19833, T19831};
  assign T19831 = $signed(T19832) / $signed(22'h100000);
  assign T19832 = $signed(30'h187de2a6) * $signed(16'hffff);
  assign T19833 = T19831[6'h2d:6'h2d];
  assign T19834 = $signed(T19835) / $signed(22'h100000);
  assign T19835 = $signed(31'h3b20d79e) * $signed(16'h0);
  assign twiddle4_1_129_imag = T19840 + T19836;
  assign T19836 = {T19839, T19837};
  assign T19837 = $signed(T19838) / $signed(22'h100000);
  assign T19838 = $signed(30'h18ac4b86) * $signed(16'hffff);
  assign T19839 = T19837[6'h2d:6'h2d];
  assign T19840 = $signed(T19841) / $signed(22'h100000);
  assign T19841 = $signed(31'h3b0d8908) * $signed(16'h0);
  assign T19842 = T18725[1'h0:1'h0];
  assign T19843 = T19856 ? twiddle4_1_131_imag : twiddle4_1_130_imag;
  assign twiddle4_1_130_imag = T19848 + T19844;
  assign T19844 = {T19847, T19845};
  assign T19845 = $signed(T19846) / $signed(22'h100000);
  assign T19846 = $signed(30'h18daa52e) * $signed(16'hffff);
  assign T19847 = T19845[6'h2d:6'h2d];
  assign T19848 = $signed(T19849) / $signed(22'h100000);
  assign T19849 = $signed(31'h3afa1605) * $signed(16'h0);
  assign twiddle4_1_131_imag = T19854 + T19850;
  assign T19850 = {T19853, T19851};
  assign T19851 = $signed(T19852) / $signed(22'h100000);
  assign T19852 = $signed(30'h1908ef81) * $signed(16'hffff);
  assign T19853 = T19851[6'h2d:6'h2d];
  assign T19854 = $signed(T19855) / $signed(22'h100000);
  assign T19855 = $signed(31'h3ae67ea1) * $signed(16'h0);
  assign T19856 = T18725[1'h0:1'h0];
  assign T19857 = T18725[1'h1:1'h1];
  assign T19858 = T19887 ? T19873 : T19859;
  assign T19859 = T19872 ? twiddle4_1_133_imag : twiddle4_1_132_imag;
  assign twiddle4_1_132_imag = T19864 + T19860;
  assign T19860 = {T19863, T19861};
  assign T19861 = $signed(T19862) / $signed(22'h100000);
  assign T19862 = $signed(30'h19372a63) * $signed(16'hffff);
  assign T19863 = T19861[6'h2d:6'h2d];
  assign T19864 = $signed(T19865) / $signed(22'h100000);
  assign T19865 = $signed(31'h3ad2c2e7) * $signed(16'h0);
  assign twiddle4_1_133_imag = T19870 + T19866;
  assign T19866 = {T19869, T19867};
  assign T19867 = $signed(T19868) / $signed(22'h100000);
  assign T19868 = $signed(30'h196555b7) * $signed(16'hffff);
  assign T19869 = T19867[6'h2d:6'h2d];
  assign T19870 = $signed(T19871) / $signed(22'h100000);
  assign T19871 = $signed(31'h3abee2e5) * $signed(16'h0);
  assign T19872 = T18725[1'h0:1'h0];
  assign T19873 = T19886 ? twiddle4_1_135_imag : twiddle4_1_134_imag;
  assign twiddle4_1_134_imag = T19878 + T19874;
  assign T19874 = {T19877, T19875};
  assign T19875 = $signed(T19876) / $signed(22'h100000);
  assign T19876 = $signed(30'h19937161) * $signed(16'hffff);
  assign T19877 = T19875[6'h2d:6'h2d];
  assign T19878 = $signed(T19879) / $signed(22'h100000);
  assign T19879 = $signed(31'h3aaadea5) * $signed(16'h0);
  assign twiddle4_1_135_imag = T19884 + T19880;
  assign T19880 = {T19883, T19881};
  assign T19881 = $signed(T19882) / $signed(22'h100000);
  assign T19882 = $signed(30'h19c17d44) * $signed(16'hffff);
  assign T19883 = T19881[6'h2d:6'h2d];
  assign T19884 = $signed(T19885) / $signed(22'h100000);
  assign T19885 = $signed(31'h3a96b636) * $signed(16'h0);
  assign T19886 = T18725[1'h0:1'h0];
  assign T19887 = T18725[1'h1:1'h1];
  assign T19888 = T18725[2'h2:2'h2];
  assign T19889 = T19950 ? T19920 : T19890;
  assign T19890 = T19919 ? T19905 : T19891;
  assign T19891 = T19904 ? twiddle4_1_137_imag : twiddle4_1_136_imag;
  assign twiddle4_1_136_imag = T19896 + T19892;
  assign T19892 = {T19895, T19893};
  assign T19893 = $signed(T19894) / $signed(22'h100000);
  assign T19894 = $signed(30'h19ef7943) * $signed(16'hffff);
  assign T19895 = T19893[6'h2d:6'h2d];
  assign T19896 = $signed(T19897) / $signed(22'h100000);
  assign T19897 = $signed(31'h3a8269a2) * $signed(16'h0);
  assign twiddle4_1_137_imag = T19902 + T19898;
  assign T19898 = {T19901, T19899};
  assign T19899 = $signed(T19900) / $signed(22'h100000);
  assign T19900 = $signed(30'h1a1d6543) * $signed(16'hffff);
  assign T19901 = T19899[6'h2d:6'h2d];
  assign T19902 = $signed(T19903) / $signed(22'h100000);
  assign T19903 = $signed(31'h3a6df8f7) * $signed(16'h0);
  assign T19904 = T18725[1'h0:1'h0];
  assign T19905 = T19918 ? twiddle4_1_139_imag : twiddle4_1_138_imag;
  assign twiddle4_1_138_imag = T19910 + T19906;
  assign T19906 = {T19909, T19907};
  assign T19907 = $signed(T19908) / $signed(22'h100000);
  assign T19908 = $signed(30'h1a4b4127) * $signed(16'hffff);
  assign T19909 = T19907[6'h2d:6'h2d];
  assign T19910 = $signed(T19911) / $signed(22'h100000);
  assign T19911 = $signed(31'h3a596441) * $signed(16'h0);
  assign twiddle4_1_139_imag = T19916 + T19912;
  assign T19912 = {T19915, T19913};
  assign T19913 = $signed(T19914) / $signed(22'h100000);
  assign T19914 = $signed(30'h1a790cd3) * $signed(16'hffff);
  assign T19915 = T19913[6'h2d:6'h2d];
  assign T19916 = $signed(T19917) / $signed(22'h100000);
  assign T19917 = $signed(31'h3a44ab8d) * $signed(16'h0);
  assign T19918 = T18725[1'h0:1'h0];
  assign T19919 = T18725[1'h1:1'h1];
  assign T19920 = T19949 ? T19935 : T19921;
  assign T19921 = T19934 ? twiddle4_1_141_imag : twiddle4_1_140_imag;
  assign twiddle4_1_140_imag = T19926 + T19922;
  assign T19922 = {T19925, T19923};
  assign T19923 = $signed(T19924) / $signed(22'h100000);
  assign T19924 = $signed(30'h1aa6c82b) * $signed(16'hffff);
  assign T19925 = T19923[6'h2d:6'h2d];
  assign T19926 = $signed(T19927) / $signed(22'h100000);
  assign T19927 = $signed(31'h3a2fcee8) * $signed(16'h0);
  assign twiddle4_1_141_imag = T19932 + T19928;
  assign T19928 = {T19931, T19929};
  assign T19929 = $signed(T19930) / $signed(22'h100000);
  assign T19930 = $signed(30'h1ad47312) * $signed(16'hffff);
  assign T19931 = T19929[6'h2d:6'h2d];
  assign T19932 = $signed(T19933) / $signed(22'h100000);
  assign T19933 = $signed(31'h3a1ace5e) * $signed(16'h0);
  assign T19934 = T18725[1'h0:1'h0];
  assign T19935 = T19948 ? twiddle4_1_143_imag : twiddle4_1_142_imag;
  assign twiddle4_1_142_imag = T19940 + T19936;
  assign T19936 = {T19939, T19937};
  assign T19937 = $signed(T19938) / $signed(22'h100000);
  assign T19938 = $signed(30'h1b020d6c) * $signed(16'hffff);
  assign T19939 = T19937[6'h2d:6'h2d];
  assign T19940 = $signed(T19941) / $signed(22'h100000);
  assign T19941 = $signed(31'h3a05a9fd) * $signed(16'h0);
  assign twiddle4_1_143_imag = T19946 + T19942;
  assign T19942 = {T19945, T19943};
  assign T19943 = $signed(T19944) / $signed(22'h100000);
  assign T19944 = $signed(30'h1b2f971d) * $signed(16'hffff);
  assign T19945 = T19943[6'h2d:6'h2d];
  assign T19946 = $signed(T19947) / $signed(22'h100000);
  assign T19947 = $signed(31'h39f061d1) * $signed(16'h0);
  assign T19948 = T18725[1'h0:1'h0];
  assign T19949 = T18725[1'h1:1'h1];
  assign T19950 = T18725[2'h2:2'h2];
  assign T19951 = T18725[2'h3:2'h3];
  assign T19952 = T20077 ? T20015 : T19953;
  assign T19953 = T20014 ? T19984 : T19954;
  assign T19954 = T19983 ? T19969 : T19955;
  assign T19955 = T19968 ? twiddle4_1_145_imag : twiddle4_1_144_imag;
  assign twiddle4_1_144_imag = T19960 + T19956;
  assign T19956 = {T19959, T19957};
  assign T19957 = $signed(T19958) / $signed(22'h100000);
  assign T19958 = $signed(30'h1b5d1009) * $signed(16'hffff);
  assign T19959 = T19957[6'h2d:6'h2d];
  assign T19960 = $signed(T19961) / $signed(22'h100000);
  assign T19961 = $signed(31'h39daf5e8) * $signed(16'h0);
  assign twiddle4_1_145_imag = T19966 + T19962;
  assign T19962 = {T19965, T19963};
  assign T19963 = $signed(T19964) / $signed(22'h100000);
  assign T19964 = $signed(30'h1b8a7814) * $signed(16'hffff);
  assign T19965 = T19963[6'h2d:6'h2d];
  assign T19966 = $signed(T19967) / $signed(22'h100000);
  assign T19967 = $signed(31'h39c5664f) * $signed(16'h0);
  assign T19968 = T18725[1'h0:1'h0];
  assign T19969 = T19982 ? twiddle4_1_147_imag : twiddle4_1_146_imag;
  assign twiddle4_1_146_imag = T19974 + T19970;
  assign T19970 = {T19973, T19971};
  assign T19971 = $signed(T19972) / $signed(22'h100000);
  assign T19972 = $signed(30'h1bb7cf23) * $signed(16'hffff);
  assign T19973 = T19971[6'h2d:6'h2d];
  assign T19974 = $signed(T19975) / $signed(22'h100000);
  assign T19975 = $signed(31'h39afb313) * $signed(16'h0);
  assign twiddle4_1_147_imag = T19980 + T19976;
  assign T19976 = {T19979, T19977};
  assign T19977 = $signed(T19978) / $signed(22'h100000);
  assign T19978 = $signed(30'h1be51517) * $signed(16'hffff);
  assign T19979 = T19977[6'h2d:6'h2d];
  assign T19980 = $signed(T19981) / $signed(22'h100000);
  assign T19981 = $signed(31'h3999dc41) * $signed(16'h0);
  assign T19982 = T18725[1'h0:1'h0];
  assign T19983 = T18725[1'h1:1'h1];
  assign T19984 = T20013 ? T19999 : T19985;
  assign T19985 = T19998 ? twiddle4_1_149_imag : twiddle4_1_148_imag;
  assign twiddle4_1_148_imag = T19990 + T19986;
  assign T19986 = {T19989, T19987};
  assign T19987 = $signed(T19988) / $signed(22'h100000);
  assign T19988 = $signed(30'h1c1249d8) * $signed(16'hffff);
  assign T19989 = T19987[6'h2d:6'h2d];
  assign T19990 = $signed(T19991) / $signed(22'h100000);
  assign T19991 = $signed(31'h3983e1e7) * $signed(16'h0);
  assign twiddle4_1_149_imag = T19996 + T19992;
  assign T19992 = {T19995, T19993};
  assign T19993 = $signed(T19994) / $signed(22'h100000);
  assign T19994 = $signed(30'h1c3f6d47) * $signed(16'hffff);
  assign T19995 = T19993[6'h2d:6'h2d];
  assign T19996 = $signed(T19997) / $signed(22'h100000);
  assign T19997 = $signed(31'h396dc414) * $signed(16'h0);
  assign T19998 = T18725[1'h0:1'h0];
  assign T19999 = T20012 ? twiddle4_1_151_imag : twiddle4_1_150_imag;
  assign twiddle4_1_150_imag = T20004 + T20000;
  assign T20000 = {T20003, T20001};
  assign T20001 = $signed(T20002) / $signed(22'h100000);
  assign T20002 = $signed(30'h1c6c7f49) * $signed(16'hffff);
  assign T20003 = T20001[6'h2d:6'h2d];
  assign T20004 = $signed(T20005) / $signed(22'h100000);
  assign T20005 = $signed(31'h395782d3) * $signed(16'h0);
  assign twiddle4_1_151_imag = T20010 + T20006;
  assign T20006 = {T20009, T20007};
  assign T20007 = $signed(T20008) / $signed(22'h100000);
  assign T20008 = $signed(30'h1c997fc3) * $signed(16'hffff);
  assign T20009 = T20007[6'h2d:6'h2d];
  assign T20010 = $signed(T20011) / $signed(22'h100000);
  assign T20011 = $signed(31'h39411e33) * $signed(16'h0);
  assign T20012 = T18725[1'h0:1'h0];
  assign T20013 = T18725[1'h1:1'h1];
  assign T20014 = T18725[2'h2:2'h2];
  assign T20015 = T20076 ? T20046 : T20016;
  assign T20016 = T20045 ? T20031 : T20017;
  assign T20017 = T20030 ? twiddle4_1_153_imag : twiddle4_1_152_imag;
  assign twiddle4_1_152_imag = T20022 + T20018;
  assign T20018 = {T20021, T20019};
  assign T20019 = $signed(T20020) / $signed(22'h100000);
  assign T20020 = $signed(30'h1cc66e99) * $signed(16'hffff);
  assign T20021 = T20019[6'h2d:6'h2d];
  assign T20022 = $signed(T20023) / $signed(22'h100000);
  assign T20023 = $signed(31'h392a9642) * $signed(16'h0);
  assign twiddle4_1_153_imag = T20028 + T20024;
  assign T20024 = {T20027, T20025};
  assign T20025 = $signed(T20026) / $signed(22'h100000);
  assign T20026 = $signed(30'h1cf34bae) * $signed(16'hffff);
  assign T20027 = T20025[6'h2d:6'h2d];
  assign T20028 = $signed(T20029) / $signed(22'h100000);
  assign T20029 = $signed(31'h3913eb0e) * $signed(16'h0);
  assign T20030 = T18725[1'h0:1'h0];
  assign T20031 = T20044 ? twiddle4_1_155_imag : twiddle4_1_154_imag;
  assign twiddle4_1_154_imag = T20036 + T20032;
  assign T20032 = {T20035, T20033};
  assign T20033 = $signed(T20034) / $signed(22'h100000);
  assign T20034 = $signed(30'h1d2016e8) * $signed(16'hffff);
  assign T20035 = T20033[6'h2d:6'h2d];
  assign T20036 = $signed(T20037) / $signed(22'h100000);
  assign T20037 = $signed(31'h38fd1ca4) * $signed(16'h0);
  assign twiddle4_1_155_imag = T20042 + T20038;
  assign T20038 = {T20041, T20039};
  assign T20039 = $signed(T20040) / $signed(22'h100000);
  assign T20040 = $signed(30'h1d4cd02b) * $signed(16'hffff);
  assign T20041 = T20039[6'h2d:6'h2d];
  assign T20042 = $signed(T20043) / $signed(22'h100000);
  assign T20043 = $signed(31'h38e62b13) * $signed(16'h0);
  assign T20044 = T18725[1'h0:1'h0];
  assign T20045 = T18725[1'h1:1'h1];
  assign T20046 = T20075 ? T20061 : T20047;
  assign T20047 = T20060 ? twiddle4_1_157_imag : twiddle4_1_156_imag;
  assign twiddle4_1_156_imag = T20052 + T20048;
  assign T20048 = {T20051, T20049};
  assign T20049 = $signed(T20050) / $signed(22'h100000);
  assign T20050 = $signed(30'h1d79775b) * $signed(16'hffff);
  assign T20051 = T20049[6'h2d:6'h2d];
  assign T20052 = $signed(T20053) / $signed(22'h100000);
  assign T20053 = $signed(31'h38cf1669) * $signed(16'h0);
  assign twiddle4_1_157_imag = T20058 + T20054;
  assign T20054 = {T20057, T20055};
  assign T20055 = $signed(T20056) / $signed(22'h100000);
  assign T20056 = $signed(30'h1da60c5c) * $signed(16'hffff);
  assign T20057 = T20055[6'h2d:6'h2d];
  assign T20058 = $signed(T20059) / $signed(22'h100000);
  assign T20059 = $signed(31'h38b7deb3) * $signed(16'h0);
  assign T20060 = T18725[1'h0:1'h0];
  assign T20061 = T20074 ? twiddle4_1_159_imag : twiddle4_1_158_imag;
  assign twiddle4_1_158_imag = T20066 + T20062;
  assign T20062 = {T20065, T20063};
  assign T20063 = $signed(T20064) / $signed(22'h100000);
  assign T20064 = $signed(30'h1dd28f14) * $signed(16'hffff);
  assign T20065 = T20063[6'h2d:6'h2d];
  assign T20066 = $signed(T20067) / $signed(22'h100000);
  assign T20067 = $signed(31'h38a08402) * $signed(16'h0);
  assign twiddle4_1_159_imag = T20072 + T20068;
  assign T20068 = {T20071, T20069};
  assign T20069 = $signed(T20070) / $signed(22'h100000);
  assign T20070 = $signed(30'h1dfeff66) * $signed(16'hffff);
  assign T20071 = T20069[6'h2d:6'h2d];
  assign T20072 = $signed(T20073) / $signed(22'h100000);
  assign T20073 = $signed(31'h38890662) * $signed(16'h0);
  assign T20074 = T18725[1'h0:1'h0];
  assign T20075 = T18725[1'h1:1'h1];
  assign T20076 = T18725[2'h2:2'h2];
  assign T20077 = T18725[2'h3:2'h3];
  assign T20078 = T18725[3'h4:3'h4];
  assign T20079 = T20290 ? T20196 : T20080;
  assign T20080 = T20195 ? T20143 : T20081;
  assign T20081 = T20142 ? T20112 : T20082;
  assign T20082 = T20111 ? T20097 : T20083;
  assign T20083 = T20096 ? twiddle4_1_161_imag : twiddle4_1_160_imag;
  assign twiddle4_1_160_imag = T20088 + T20084;
  assign T20084 = {T20087, T20085};
  assign T20085 = $signed(T20086) / $signed(22'h100000);
  assign T20086 = $signed(30'h1e2b5d38) * $signed(16'hffff);
  assign T20087 = T20085[6'h2d:6'h2d];
  assign T20088 = $signed(T20089) / $signed(22'h100000);
  assign T20089 = $signed(31'h387165e3) * $signed(16'h0);
  assign twiddle4_1_161_imag = T20094 + T20090;
  assign T20090 = {T20093, T20091};
  assign T20091 = $signed(T20092) / $signed(22'h100000);
  assign T20092 = $signed(30'h1e57a86d) * $signed(16'hffff);
  assign T20093 = T20091[6'h2d:6'h2d];
  assign T20094 = $signed(T20095) / $signed(22'h100000);
  assign T20095 = $signed(31'h3859a292) * $signed(16'h0);
  assign T20096 = T18725[1'h0:1'h0];
  assign T20097 = T20110 ? twiddle4_1_163_imag : twiddle4_1_162_imag;
  assign twiddle4_1_162_imag = T20102 + T20098;
  assign T20098 = {T20101, T20099};
  assign T20099 = $signed(T20100) / $signed(22'h100000);
  assign T20100 = $signed(30'h1e83e0ea) * $signed(16'hffff);
  assign T20101 = T20099[6'h2d:6'h2d];
  assign T20102 = $signed(T20103) / $signed(22'h100000);
  assign T20103 = $signed(31'h3841bc7f) * $signed(16'h0);
  assign twiddle4_1_163_imag = T20108 + T20104;
  assign T20104 = {T20107, T20105};
  assign T20105 = $signed(T20106) / $signed(22'h100000);
  assign T20106 = $signed(30'h1eb00695) * $signed(16'hffff);
  assign T20107 = T20105[6'h2d:6'h2d];
  assign T20108 = $signed(T20109) / $signed(22'h100000);
  assign T20109 = $signed(31'h3829b3b8) * $signed(16'h0);
  assign T20110 = T18725[1'h0:1'h0];
  assign T20111 = T18725[1'h1:1'h1];
  assign T20112 = T20141 ? T20127 : T20113;
  assign T20113 = T20126 ? twiddle4_1_165_imag : twiddle4_1_164_imag;
  assign twiddle4_1_164_imag = T20118 + T20114;
  assign T20114 = {T20117, T20115};
  assign T20115 = $signed(T20116) / $signed(22'h100000);
  assign T20116 = $signed(30'h1edc1952) * $signed(16'hffff);
  assign T20117 = T20115[6'h2d:6'h2d];
  assign T20118 = $signed(T20119) / $signed(22'h100000);
  assign T20119 = $signed(31'h3811884c) * $signed(16'h0);
  assign twiddle4_1_165_imag = T20124 + T20120;
  assign T20120 = {T20123, T20121};
  assign T20121 = $signed(T20122) / $signed(22'h100000);
  assign T20122 = $signed(30'h1f081906) * $signed(16'hffff);
  assign T20123 = T20121[6'h2d:6'h2d];
  assign T20124 = $signed(T20125) / $signed(22'h100000);
  assign T20125 = $signed(31'h37f93a4b) * $signed(16'h0);
  assign T20126 = T18725[1'h0:1'h0];
  assign T20127 = T20140 ? twiddle4_1_167_imag : twiddle4_1_166_imag;
  assign twiddle4_1_166_imag = T20132 + T20128;
  assign T20128 = {T20131, T20129};
  assign T20129 = $signed(T20130) / $signed(22'h100000);
  assign T20130 = $signed(30'h1f340596) * $signed(16'hffff);
  assign T20131 = T20129[6'h2d:6'h2d];
  assign T20132 = $signed(T20133) / $signed(22'h100000);
  assign T20133 = $signed(31'h37e0c9c2) * $signed(16'h0);
  assign twiddle4_1_167_imag = T20138 + T20134;
  assign T20134 = {T20137, T20135};
  assign T20135 = $signed(T20136) / $signed(22'h100000);
  assign T20136 = $signed(30'h1f5fdee6) * $signed(16'hffff);
  assign T20137 = T20135[6'h2d:6'h2d];
  assign T20138 = $signed(T20139) / $signed(22'h100000);
  assign T20139 = $signed(31'h37c836c2) * $signed(16'h0);
  assign T20140 = T18725[1'h0:1'h0];
  assign T20141 = T18725[1'h1:1'h1];
  assign T20142 = T18725[2'h2:2'h2];
  assign T20143 = T20194 ? T20172 : T20144;
  assign T20144 = T20171 ? T20159 : T20145;
  assign T20145 = T20158 ? twiddle4_1_169_imag : twiddle4_1_168_imag;
  assign twiddle4_1_168_imag = T20150 + T20146;
  assign T20146 = {T20149, T20147};
  assign T20147 = $signed(T20148) / $signed(22'h100000);
  assign T20148 = $signed(30'h1f8ba4db) * $signed(16'hffff);
  assign T20149 = T20147[6'h2d:6'h2d];
  assign T20150 = $signed(T20151) / $signed(22'h100000);
  assign T20151 = $signed(31'h37af8158) * $signed(16'h0);
  assign twiddle4_1_169_imag = T20156 + T20152;
  assign T20152 = {T20155, T20153};
  assign T20153 = $signed(T20154) / $signed(22'h100000);
  assign T20154 = $signed(30'h1fb7575c) * $signed(16'hffff);
  assign T20155 = T20153[6'h2d:6'h2d];
  assign T20156 = $signed(T20157) / $signed(22'h100000);
  assign T20157 = $signed(31'h3796a996) * $signed(16'h0);
  assign T20158 = T18725[1'h0:1'h0];
  assign T20159 = T20170 ? twiddle4_1_171_imag : twiddle4_1_170_imag;
  assign twiddle4_1_170_imag = T20164 + T20160;
  assign T20160 = {T20163, T20161};
  assign T20161 = $signed(T20162) / $signed(22'h100000);
  assign T20162 = $signed(30'h1fe2f64b) * $signed(16'hffff);
  assign T20163 = T20161[6'h2d:6'h2d];
  assign T20164 = $signed(T20165) / $signed(22'h100000);
  assign T20165 = $signed(31'h377daf89) * $signed(16'h0);
  assign twiddle4_1_171_imag = T20168 + T20166;
  assign T20166 = $signed(T20167) / $signed(22'h100000);
  assign T20167 = $signed(31'h200e8190) * $signed(16'hffff);
  assign T20168 = $signed(T20169) / $signed(22'h100000);
  assign T20169 = $signed(31'h37649341) * $signed(16'h0);
  assign T20170 = T18725[1'h0:1'h0];
  assign T20171 = T18725[1'h1:1'h1];
  assign T20172 = T20193 ? T20183 : T20173;
  assign T20173 = T20182 ? twiddle4_1_173_imag : twiddle4_1_172_imag;
  assign twiddle4_1_172_imag = T20176 + T20174;
  assign T20174 = $signed(T20175) / $signed(22'h100000);
  assign T20175 = $signed(31'h2039f90e) * $signed(16'hffff);
  assign T20176 = $signed(T20177) / $signed(22'h100000);
  assign T20177 = $signed(31'h374b54ce) * $signed(16'h0);
  assign twiddle4_1_173_imag = T20180 + T20178;
  assign T20178 = $signed(T20179) / $signed(22'h100000);
  assign T20179 = $signed(31'h20655cab) * $signed(16'hffff);
  assign T20180 = $signed(T20181) / $signed(22'h100000);
  assign T20181 = $signed(31'h3731f43f) * $signed(16'h0);
  assign T20182 = T18725[1'h0:1'h0];
  assign T20183 = T20192 ? twiddle4_1_175_imag : twiddle4_1_174_imag;
  assign twiddle4_1_174_imag = T20186 + T20184;
  assign T20184 = $signed(T20185) / $signed(22'h100000);
  assign T20185 = $signed(31'h2090ac4d) * $signed(16'hffff);
  assign T20186 = $signed(T20187) / $signed(22'h100000);
  assign T20187 = $signed(31'h371871a4) * $signed(16'h0);
  assign twiddle4_1_175_imag = T20190 + T20188;
  assign T20188 = $signed(T20189) / $signed(22'h100000);
  assign T20189 = $signed(31'h20bbe7d8) * $signed(16'hffff);
  assign T20190 = $signed(T20191) / $signed(22'h100000);
  assign T20191 = $signed(31'h36fecd0d) * $signed(16'h0);
  assign T20192 = T18725[1'h0:1'h0];
  assign T20193 = T18725[1'h1:1'h1];
  assign T20194 = T18725[2'h2:2'h2];
  assign T20195 = T18725[2'h3:2'h3];
  assign T20196 = T20289 ? T20243 : T20197;
  assign T20197 = T20242 ? T20220 : T20198;
  assign T20198 = T20219 ? T20209 : T20199;
  assign T20199 = T20208 ? twiddle4_1_177_imag : twiddle4_1_176_imag;
  assign twiddle4_1_176_imag = T20202 + T20200;
  assign T20200 = $signed(T20201) / $signed(22'h100000);
  assign T20201 = $signed(31'h20e70f32) * $signed(16'hffff);
  assign T20202 = $signed(T20203) / $signed(22'h100000);
  assign T20203 = $signed(31'h36e5068a) * $signed(16'h0);
  assign twiddle4_1_177_imag = T20206 + T20204;
  assign T20204 = $signed(T20205) / $signed(22'h100000);
  assign T20205 = $signed(31'h21122240) * $signed(16'hffff);
  assign T20206 = $signed(T20207) / $signed(22'h100000);
  assign T20207 = $signed(31'h36cb1e29) * $signed(16'h0);
  assign T20208 = T18725[1'h0:1'h0];
  assign T20209 = T20218 ? twiddle4_1_179_imag : twiddle4_1_178_imag;
  assign twiddle4_1_178_imag = T20212 + T20210;
  assign T20210 = $signed(T20211) / $signed(22'h100000);
  assign T20211 = $signed(31'h213d20e8) * $signed(16'hffff);
  assign T20212 = $signed(T20213) / $signed(22'h100000);
  assign T20213 = $signed(31'h36b113fd) * $signed(16'h0);
  assign twiddle4_1_179_imag = T20216 + T20214;
  assign T20214 = $signed(T20215) / $signed(22'h100000);
  assign T20215 = $signed(31'h21680b0f) * $signed(16'hffff);
  assign T20216 = $signed(T20217) / $signed(22'h100000);
  assign T20217 = $signed(31'h3696e813) * $signed(16'h0);
  assign T20218 = T18725[1'h0:1'h0];
  assign T20219 = T18725[1'h1:1'h1];
  assign T20220 = T20241 ? T20231 : T20221;
  assign T20221 = T20230 ? twiddle4_1_181_imag : twiddle4_1_180_imag;
  assign twiddle4_1_180_imag = T20224 + T20222;
  assign T20222 = $signed(T20223) / $signed(22'h100000);
  assign T20223 = $signed(31'h2192e09a) * $signed(16'hffff);
  assign T20224 = $signed(T20225) / $signed(22'h100000);
  assign T20225 = $signed(31'h367c9a7d) * $signed(16'h0);
  assign twiddle4_1_181_imag = T20228 + T20226;
  assign T20226 = $signed(T20227) / $signed(22'h100000);
  assign T20227 = $signed(31'h21bda170) * $signed(16'hffff);
  assign T20228 = $signed(T20229) / $signed(22'h100000);
  assign T20229 = $signed(31'h36622b4b) * $signed(16'h0);
  assign T20230 = T18725[1'h0:1'h0];
  assign T20231 = T20240 ? twiddle4_1_183_imag : twiddle4_1_182_imag;
  assign twiddle4_1_182_imag = T20234 + T20232;
  assign T20232 = $signed(T20233) / $signed(22'h100000);
  assign T20233 = $signed(31'h21e84d76) * $signed(16'hffff);
  assign T20234 = $signed(T20235) / $signed(22'h100000);
  assign T20235 = $signed(31'h36479a8e) * $signed(16'h0);
  assign twiddle4_1_183_imag = T20238 + T20236;
  assign T20236 = $signed(T20237) / $signed(22'h100000);
  assign T20237 = $signed(31'h2212e491) * $signed(16'hffff);
  assign T20238 = $signed(T20239) / $signed(22'h100000);
  assign T20239 = $signed(31'h362ce854) * $signed(16'h0);
  assign T20240 = T18725[1'h0:1'h0];
  assign T20241 = T18725[1'h1:1'h1];
  assign T20242 = T18725[2'h2:2'h2];
  assign T20243 = T20288 ? T20266 : T20244;
  assign T20244 = T20265 ? T20255 : T20245;
  assign T20245 = T20254 ? twiddle4_1_185_imag : twiddle4_1_184_imag;
  assign twiddle4_1_184_imag = T20248 + T20246;
  assign T20246 = $signed(T20247) / $signed(22'h100000);
  assign T20247 = $signed(31'h223d66a8) * $signed(16'hffff);
  assign T20248 = $signed(T20249) / $signed(22'h100000);
  assign T20249 = $signed(31'h361214b0) * $signed(16'h0);
  assign twiddle4_1_185_imag = T20252 + T20250;
  assign T20250 = $signed(T20251) / $signed(22'h100000);
  assign T20251 = $signed(31'h2267d39f) * $signed(16'hffff);
  assign T20252 = $signed(T20253) / $signed(22'h100000);
  assign T20253 = $signed(31'h35f71fb1) * $signed(16'h0);
  assign T20254 = T18725[1'h0:1'h0];
  assign T20255 = T20264 ? twiddle4_1_187_imag : twiddle4_1_186_imag;
  assign twiddle4_1_186_imag = T20258 + T20256;
  assign T20256 = $signed(T20257) / $signed(22'h100000);
  assign T20257 = $signed(31'h22922b5e) * $signed(16'hffff);
  assign T20258 = $signed(T20259) / $signed(22'h100000);
  assign T20259 = $signed(31'h35dc0968) * $signed(16'h0);
  assign twiddle4_1_187_imag = T20262 + T20260;
  assign T20260 = $signed(T20261) / $signed(22'h100000);
  assign T20261 = $signed(31'h22bc6dc9) * $signed(16'hffff);
  assign T20262 = $signed(T20263) / $signed(22'h100000);
  assign T20263 = $signed(31'h35c0d1e6) * $signed(16'h0);
  assign T20264 = T18725[1'h0:1'h0];
  assign T20265 = T18725[1'h1:1'h1];
  assign T20266 = T20287 ? T20277 : T20267;
  assign T20267 = T20276 ? twiddle4_1_189_imag : twiddle4_1_188_imag;
  assign twiddle4_1_188_imag = T20270 + T20268;
  assign T20268 = $signed(T20269) / $signed(22'h100000);
  assign T20269 = $signed(31'h22e69ac7) * $signed(16'hffff);
  assign T20270 = $signed(T20271) / $signed(22'h100000);
  assign T20271 = $signed(31'h35a5793c) * $signed(16'h0);
  assign twiddle4_1_189_imag = T20274 + T20272;
  assign T20272 = $signed(T20273) / $signed(22'h100000);
  assign T20273 = $signed(31'h2310b23e) * $signed(16'hffff);
  assign T20274 = $signed(T20275) / $signed(22'h100000);
  assign T20275 = $signed(31'h3589ff7a) * $signed(16'h0);
  assign T20276 = T18725[1'h0:1'h0];
  assign T20277 = T20286 ? twiddle4_1_191_imag : twiddle4_1_190_imag;
  assign twiddle4_1_190_imag = T20280 + T20278;
  assign T20278 = $signed(T20279) / $signed(22'h100000);
  assign T20279 = $signed(31'h233ab413) * $signed(16'hffff);
  assign T20280 = $signed(T20281) / $signed(22'h100000);
  assign T20281 = $signed(31'h356e64b2) * $signed(16'h0);
  assign twiddle4_1_191_imag = T20284 + T20282;
  assign T20282 = $signed(T20283) / $signed(22'h100000);
  assign T20283 = $signed(31'h2364a02e) * $signed(16'hffff);
  assign T20284 = $signed(T20285) / $signed(22'h100000);
  assign T20285 = $signed(31'h3552a8f4) * $signed(16'h0);
  assign T20286 = T18725[1'h0:1'h0];
  assign T20287 = T18725[1'h1:1'h1];
  assign T20288 = T18725[2'h2:2'h2];
  assign T20289 = T18725[2'h3:2'h3];
  assign T20290 = T18725[3'h4:3'h4];
  assign T20291 = T18725[3'h5:3'h5];
  assign T20292 = T20673 ? T20483 : T20293;
  assign T20293 = T20482 ? T20388 : T20294;
  assign T20294 = T20387 ? T20341 : T20295;
  assign T20295 = T20340 ? T20318 : T20296;
  assign T20296 = T20317 ? T20307 : T20297;
  assign T20297 = T20306 ? twiddle4_1_193_imag : twiddle4_1_192_imag;
  assign twiddle4_1_192_imag = T20300 + T20298;
  assign T20298 = $signed(T20299) / $signed(22'h100000);
  assign T20299 = $signed(31'h238e7673) * $signed(16'hffff);
  assign T20300 = $signed(T20301) / $signed(22'h100000);
  assign T20301 = $signed(31'h3536cc52) * $signed(16'h0);
  assign twiddle4_1_193_imag = T20304 + T20302;
  assign T20302 = $signed(T20303) / $signed(22'h100000);
  assign T20303 = $signed(31'h23b836c9) * $signed(16'hffff);
  assign T20304 = $signed(T20305) / $signed(22'h100000);
  assign T20305 = $signed(31'h351acedc) * $signed(16'h0);
  assign T20306 = T18725[1'h0:1'h0];
  assign T20307 = T20316 ? twiddle4_1_195_imag : twiddle4_1_194_imag;
  assign twiddle4_1_194_imag = T20310 + T20308;
  assign T20308 = $signed(T20309) / $signed(22'h100000);
  assign T20309 = $signed(31'h23e1e117) * $signed(16'hffff);
  assign T20310 = $signed(T20311) / $signed(22'h100000);
  assign T20311 = $signed(31'h34feb0a5) * $signed(16'h0);
  assign twiddle4_1_195_imag = T20314 + T20312;
  assign T20312 = $signed(T20313) / $signed(22'h100000);
  assign T20313 = $signed(31'h240b7542) * $signed(16'hffff);
  assign T20314 = $signed(T20315) / $signed(22'h100000);
  assign T20315 = $signed(31'h34e271bd) * $signed(16'h0);
  assign T20316 = T18725[1'h0:1'h0];
  assign T20317 = T18725[1'h1:1'h1];
  assign T20318 = T20339 ? T20329 : T20319;
  assign T20319 = T20328 ? twiddle4_1_197_imag : twiddle4_1_196_imag;
  assign twiddle4_1_196_imag = T20322 + T20320;
  assign T20320 = $signed(T20321) / $signed(22'h100000);
  assign T20321 = $signed(31'h2434f332) * $signed(16'hffff);
  assign T20322 = $signed(T20323) / $signed(22'h100000);
  assign T20323 = $signed(31'h34c61236) * $signed(16'h0);
  assign twiddle4_1_197_imag = T20326 + T20324;
  assign T20324 = $signed(T20325) / $signed(22'h100000);
  assign T20325 = $signed(31'h245e5acc) * $signed(16'hffff);
  assign T20326 = $signed(T20327) / $signed(22'h100000);
  assign T20327 = $signed(31'h34a99221) * $signed(16'h0);
  assign T20328 = T18725[1'h0:1'h0];
  assign T20329 = T20338 ? twiddle4_1_199_imag : twiddle4_1_198_imag;
  assign twiddle4_1_198_imag = T20332 + T20330;
  assign T20330 = $signed(T20331) / $signed(22'h100000);
  assign T20331 = $signed(31'h2487abf7) * $signed(16'hffff);
  assign T20332 = $signed(T20333) / $signed(22'h100000);
  assign T20333 = $signed(31'h348cf190) * $signed(16'h0);
  assign twiddle4_1_199_imag = T20336 + T20334;
  assign T20334 = $signed(T20335) / $signed(22'h100000);
  assign T20335 = $signed(31'h24b0e699) * $signed(16'hffff);
  assign T20336 = $signed(T20337) / $signed(22'h100000);
  assign T20337 = $signed(31'h34703094) * $signed(16'h0);
  assign T20338 = T18725[1'h0:1'h0];
  assign T20339 = T18725[1'h1:1'h1];
  assign T20340 = T18725[2'h2:2'h2];
  assign T20341 = T20386 ? T20364 : T20342;
  assign T20342 = T20363 ? T20353 : T20343;
  assign T20343 = T20352 ? twiddle4_1_201_imag : twiddle4_1_200_imag;
  assign twiddle4_1_200_imag = T20346 + T20344;
  assign T20344 = $signed(T20345) / $signed(22'h100000);
  assign T20345 = $signed(31'h24da0a99) * $signed(16'hffff);
  assign T20346 = $signed(T20347) / $signed(22'h100000);
  assign T20347 = $signed(31'h34534f40) * $signed(16'h0);
  assign twiddle4_1_201_imag = T20350 + T20348;
  assign T20348 = $signed(T20349) / $signed(22'h100000);
  assign T20349 = $signed(31'h250317de) * $signed(16'hffff);
  assign T20350 = $signed(T20351) / $signed(22'h100000);
  assign T20351 = $signed(31'h34364da5) * $signed(16'h0);
  assign T20352 = T18725[1'h0:1'h0];
  assign T20353 = T20362 ? twiddle4_1_203_imag : twiddle4_1_202_imag;
  assign twiddle4_1_202_imag = T20356 + T20354;
  assign T20354 = $signed(T20355) / $signed(22'h100000);
  assign T20355 = $signed(31'h252c0e4e) * $signed(16'hffff);
  assign T20356 = $signed(T20357) / $signed(22'h100000);
  assign T20357 = $signed(31'h34192bd5) * $signed(16'h0);
  assign twiddle4_1_203_imag = T20360 + T20358;
  assign T20358 = $signed(T20359) / $signed(22'h100000);
  assign T20359 = $signed(31'h2554edd0) * $signed(16'hffff);
  assign T20360 = $signed(T20361) / $signed(22'h100000);
  assign T20361 = $signed(31'h33fbe9e2) * $signed(16'h0);
  assign T20362 = T18725[1'h0:1'h0];
  assign T20363 = T18725[1'h1:1'h1];
  assign T20364 = T20385 ? T20375 : T20365;
  assign T20365 = T20374 ? twiddle4_1_205_imag : twiddle4_1_204_imag;
  assign twiddle4_1_204_imag = T20368 + T20366;
  assign T20366 = $signed(T20367) / $signed(22'h100000);
  assign T20367 = $signed(31'h257db64b) * $signed(16'hffff);
  assign T20368 = $signed(T20369) / $signed(22'h100000);
  assign T20369 = $signed(31'h33de87de) * $signed(16'h0);
  assign twiddle4_1_205_imag = T20372 + T20370;
  assign T20370 = $signed(T20371) / $signed(22'h100000);
  assign T20371 = $signed(31'h25a667a6) * $signed(16'hffff);
  assign T20372 = $signed(T20373) / $signed(22'h100000);
  assign T20373 = $signed(31'h33c105db) * $signed(16'h0);
  assign T20374 = T18725[1'h0:1'h0];
  assign T20375 = T20384 ? twiddle4_1_207_imag : twiddle4_1_206_imag;
  assign twiddle4_1_206_imag = T20378 + T20376;
  assign T20376 = $signed(T20377) / $signed(22'h100000);
  assign T20377 = $signed(31'h25cf01c7) * $signed(16'hffff);
  assign T20378 = $signed(T20379) / $signed(22'h100000);
  assign T20379 = $signed(31'h33a363eb) * $signed(16'h0);
  assign twiddle4_1_207_imag = T20382 + T20380;
  assign T20380 = $signed(T20381) / $signed(22'h100000);
  assign T20381 = $signed(31'h25f78496) * $signed(16'hffff);
  assign T20382 = $signed(T20383) / $signed(22'h100000);
  assign T20383 = $signed(31'h3385a221) * $signed(16'h0);
  assign T20384 = T18725[1'h0:1'h0];
  assign T20385 = T18725[1'h1:1'h1];
  assign T20386 = T18725[2'h2:2'h2];
  assign T20387 = T18725[2'h3:2'h3];
  assign T20388 = T20481 ? T20435 : T20389;
  assign T20389 = T20434 ? T20412 : T20390;
  assign T20390 = T20411 ? T20401 : T20391;
  assign T20391 = T20400 ? twiddle4_1_209_imag : twiddle4_1_208_imag;
  assign twiddle4_1_208_imag = T20394 + T20392;
  assign T20392 = $signed(T20393) / $signed(22'h100000);
  assign T20393 = $signed(31'h261feff9) * $signed(16'hffff);
  assign T20394 = $signed(T20395) / $signed(22'h100000);
  assign T20395 = $signed(31'h3367c08f) * $signed(16'h0);
  assign twiddle4_1_209_imag = T20398 + T20396;
  assign T20396 = $signed(T20397) / $signed(22'h100000);
  assign T20397 = $signed(31'h264843d8) * $signed(16'hffff);
  assign T20398 = $signed(T20399) / $signed(22'h100000);
  assign T20399 = $signed(31'h3349bf48) * $signed(16'h0);
  assign T20400 = T18725[1'h0:1'h0];
  assign T20401 = T20410 ? twiddle4_1_211_imag : twiddle4_1_210_imag;
  assign twiddle4_1_210_imag = T20404 + T20402;
  assign T20402 = $signed(T20403) / $signed(22'h100000);
  assign T20403 = $signed(31'h2670801a) * $signed(16'hffff);
  assign T20404 = $signed(T20405) / $signed(22'h100000);
  assign T20405 = $signed(31'h332b9e5d) * $signed(16'h0);
  assign twiddle4_1_211_imag = T20408 + T20406;
  assign T20406 = $signed(T20407) / $signed(22'h100000);
  assign T20407 = $signed(31'h2698a4a5) * $signed(16'hffff);
  assign T20408 = $signed(T20409) / $signed(22'h100000);
  assign T20409 = $signed(31'h330d5de2) * $signed(16'h0);
  assign T20410 = T18725[1'h0:1'h0];
  assign T20411 = T18725[1'h1:1'h1];
  assign T20412 = T20433 ? T20423 : T20413;
  assign T20413 = T20422 ? twiddle4_1_213_imag : twiddle4_1_212_imag;
  assign twiddle4_1_212_imag = T20416 + T20414;
  assign T20414 = $signed(T20415) / $signed(22'h100000);
  assign T20415 = $signed(31'h26c0b162) * $signed(16'hffff);
  assign T20416 = $signed(T20417) / $signed(22'h100000);
  assign T20417 = $signed(31'h32eefde9) * $signed(16'h0);
  assign twiddle4_1_213_imag = T20420 + T20418;
  assign T20418 = $signed(T20419) / $signed(22'h100000);
  assign T20419 = $signed(31'h26e8a637) * $signed(16'hffff);
  assign T20420 = $signed(T20421) / $signed(22'h100000);
  assign T20421 = $signed(31'h32d07e85) * $signed(16'h0);
  assign T20422 = T18725[1'h0:1'h0];
  assign T20423 = T20432 ? twiddle4_1_215_imag : twiddle4_1_214_imag;
  assign twiddle4_1_214_imag = T20426 + T20424;
  assign T20424 = $signed(T20425) / $signed(22'h100000);
  assign T20425 = $signed(31'h2710830b) * $signed(16'hffff);
  assign T20426 = $signed(T20427) / $signed(22'h100000);
  assign T20427 = $signed(31'h32b1dfc9) * $signed(16'h0);
  assign twiddle4_1_215_imag = T20430 + T20428;
  assign T20428 = $signed(T20429) / $signed(22'h100000);
  assign T20429 = $signed(31'h273847c7) * $signed(16'hffff);
  assign T20430 = $signed(T20431) / $signed(22'h100000);
  assign T20431 = $signed(31'h329321c7) * $signed(16'h0);
  assign T20432 = T18725[1'h0:1'h0];
  assign T20433 = T18725[1'h1:1'h1];
  assign T20434 = T18725[2'h2:2'h2];
  assign T20435 = T20480 ? T20458 : T20436;
  assign T20436 = T20457 ? T20447 : T20437;
  assign T20437 = T20446 ? twiddle4_1_217_imag : twiddle4_1_216_imag;
  assign twiddle4_1_216_imag = T20440 + T20438;
  assign T20438 = $signed(T20439) / $signed(22'h100000);
  assign T20439 = $signed(31'h275ff452) * $signed(16'hffff);
  assign T20440 = $signed(T20441) / $signed(22'h100000);
  assign T20441 = $signed(31'h32744493) * $signed(16'h0);
  assign twiddle4_1_217_imag = T20444 + T20442;
  assign T20442 = $signed(T20443) / $signed(22'h100000);
  assign T20443 = $signed(31'h27878893) * $signed(16'hffff);
  assign T20444 = $signed(T20445) / $signed(22'h100000);
  assign T20445 = $signed(31'h3255483f) * $signed(16'h0);
  assign T20446 = T18725[1'h0:1'h0];
  assign T20447 = T20456 ? twiddle4_1_219_imag : twiddle4_1_218_imag;
  assign twiddle4_1_218_imag = T20450 + T20448;
  assign T20448 = $signed(T20449) / $signed(22'h100000);
  assign T20449 = $signed(31'h27af0471) * $signed(16'hffff);
  assign T20450 = $signed(T20451) / $signed(22'h100000);
  assign T20451 = $signed(31'h32362cdf) * $signed(16'h0);
  assign twiddle4_1_219_imag = T20454 + T20452;
  assign T20452 = $signed(T20453) / $signed(22'h100000);
  assign T20453 = $signed(31'h27d667d5) * $signed(16'hffff);
  assign T20454 = $signed(T20455) / $signed(22'h100000);
  assign T20455 = $signed(31'h3216f286) * $signed(16'h0);
  assign T20456 = T18725[1'h0:1'h0];
  assign T20457 = T18725[1'h1:1'h1];
  assign T20458 = T20479 ? T20469 : T20459;
  assign T20459 = T20468 ? twiddle4_1_221_imag : twiddle4_1_220_imag;
  assign twiddle4_1_220_imag = T20462 + T20460;
  assign T20460 = $signed(T20461) / $signed(22'h100000);
  assign T20461 = $signed(31'h27fdb2a6) * $signed(16'hffff);
  assign T20462 = $signed(T20463) / $signed(22'h100000);
  assign T20463 = $signed(31'h31f79947) * $signed(16'h0);
  assign twiddle4_1_221_imag = T20466 + T20464;
  assign T20464 = $signed(T20465) / $signed(22'h100000);
  assign T20465 = $signed(31'h2824e4cc) * $signed(16'hffff);
  assign T20466 = $signed(T20467) / $signed(22'h100000);
  assign T20467 = $signed(31'h31d82136) * $signed(16'h0);
  assign T20468 = T18725[1'h0:1'h0];
  assign T20469 = T20478 ? twiddle4_1_223_imag : twiddle4_1_222_imag;
  assign twiddle4_1_222_imag = T20472 + T20470;
  assign T20470 = $signed(T20471) / $signed(22'h100000);
  assign T20471 = $signed(31'h284bfe2f) * $signed(16'hffff);
  assign T20472 = $signed(T20473) / $signed(22'h100000);
  assign T20473 = $signed(31'h31b88a66) * $signed(16'h0);
  assign twiddle4_1_223_imag = T20476 + T20474;
  assign T20474 = $signed(T20475) / $signed(22'h100000);
  assign T20475 = $signed(31'h2872feb6) * $signed(16'hffff);
  assign T20476 = $signed(T20477) / $signed(22'h100000);
  assign T20477 = $signed(31'h3198d4ea) * $signed(16'h0);
  assign T20478 = T18725[1'h0:1'h0];
  assign T20479 = T18725[1'h1:1'h1];
  assign T20480 = T18725[2'h2:2'h2];
  assign T20481 = T18725[2'h3:2'h3];
  assign T20482 = T18725[3'h4:3'h4];
  assign T20483 = T20672 ? T20578 : T20484;
  assign T20484 = T20577 ? T20531 : T20485;
  assign T20485 = T20530 ? T20508 : T20486;
  assign T20486 = T20507 ? T20497 : T20487;
  assign T20487 = T20496 ? twiddle4_1_225_imag : twiddle4_1_224_imag;
  assign twiddle4_1_224_imag = T20490 + T20488;
  assign T20488 = $signed(T20489) / $signed(22'h100000);
  assign T20489 = $signed(31'h2899e64a) * $signed(16'hffff);
  assign T20490 = $signed(T20491) / $signed(22'h100000);
  assign T20491 = $signed(31'h317900d6) * $signed(16'h0);
  assign twiddle4_1_225_imag = T20494 + T20492;
  assign T20492 = $signed(T20493) / $signed(22'h100000);
  assign T20493 = $signed(31'h28c0b4d2) * $signed(16'hffff);
  assign T20494 = $signed(T20495) / $signed(22'h100000);
  assign T20495 = $signed(31'h31590e3d) * $signed(16'h0);
  assign T20496 = T18725[1'h0:1'h0];
  assign T20497 = T20506 ? twiddle4_1_227_imag : twiddle4_1_226_imag;
  assign twiddle4_1_226_imag = T20500 + T20498;
  assign T20498 = $signed(T20499) / $signed(22'h100000);
  assign T20499 = $signed(31'h28e76a37) * $signed(16'hffff);
  assign T20500 = $signed(T20501) / $signed(22'h100000);
  assign T20501 = $signed(31'h3138fd34) * $signed(16'h0);
  assign twiddle4_1_227_imag = T20504 + T20502;
  assign T20502 = $signed(T20503) / $signed(22'h100000);
  assign T20503 = $signed(31'h290e0660) * $signed(16'hffff);
  assign T20504 = $signed(T20505) / $signed(22'h100000);
  assign T20505 = $signed(31'h3118cdce) * $signed(16'h0);
  assign T20506 = T18725[1'h0:1'h0];
  assign T20507 = T18725[1'h1:1'h1];
  assign T20508 = T20529 ? T20519 : T20509;
  assign T20509 = T20518 ? twiddle4_1_229_imag : twiddle4_1_228_imag;
  assign twiddle4_1_228_imag = T20512 + T20510;
  assign T20510 = $signed(T20511) / $signed(22'h100000);
  assign T20511 = $signed(31'h29348937) * $signed(16'hffff);
  assign T20512 = $signed(T20513) / $signed(22'h100000);
  assign T20513 = $signed(31'h30f8801f) * $signed(16'h0);
  assign twiddle4_1_229_imag = T20516 + T20514;
  assign T20514 = $signed(T20515) / $signed(22'h100000);
  assign T20515 = $signed(31'h295af2a2) * $signed(16'hffff);
  assign T20516 = $signed(T20517) / $signed(22'h100000);
  assign T20517 = $signed(31'h30d8143b) * $signed(16'h0);
  assign T20518 = T18725[1'h0:1'h0];
  assign T20519 = T20528 ? twiddle4_1_231_imag : twiddle4_1_230_imag;
  assign twiddle4_1_230_imag = T20522 + T20520;
  assign T20520 = $signed(T20521) / $signed(22'h100000);
  assign T20521 = $signed(31'h2981428b) * $signed(16'hffff);
  assign T20522 = $signed(T20523) / $signed(22'h100000);
  assign T20523 = $signed(31'h30b78a35) * $signed(16'h0);
  assign twiddle4_1_231_imag = T20526 + T20524;
  assign T20524 = $signed(T20525) / $signed(22'h100000);
  assign T20525 = $signed(31'h29a778da) * $signed(16'hffff);
  assign T20526 = $signed(T20527) / $signed(22'h100000);
  assign T20527 = $signed(31'h3096e223) * $signed(16'h0);
  assign T20528 = T18725[1'h0:1'h0];
  assign T20529 = T18725[1'h1:1'h1];
  assign T20530 = T18725[2'h2:2'h2];
  assign T20531 = T20576 ? T20554 : T20532;
  assign T20532 = T20553 ? T20543 : T20533;
  assign T20533 = T20542 ? twiddle4_1_233_imag : twiddle4_1_232_imag;
  assign twiddle4_1_232_imag = T20536 + T20534;
  assign T20534 = $signed(T20535) / $signed(22'h100000);
  assign T20535 = $signed(31'h29cd9577) * $signed(16'hffff);
  assign T20536 = $signed(T20537) / $signed(22'h100000);
  assign T20537 = $signed(31'h30761c17) * $signed(16'h0);
  assign twiddle4_1_233_imag = T20540 + T20538;
  assign T20538 = $signed(T20539) / $signed(22'h100000);
  assign T20539 = $signed(31'h29f3984b) * $signed(16'hffff);
  assign T20540 = $signed(T20541) / $signed(22'h100000);
  assign T20541 = $signed(31'h30553827) * $signed(16'h0);
  assign T20542 = T18725[1'h0:1'h0];
  assign T20543 = T20552 ? twiddle4_1_235_imag : twiddle4_1_234_imag;
  assign twiddle4_1_234_imag = T20546 + T20544;
  assign T20544 = $signed(T20545) / $signed(22'h100000);
  assign T20545 = $signed(31'h2a19813e) * $signed(16'hffff);
  assign T20546 = $signed(T20547) / $signed(22'h100000);
  assign T20547 = $signed(31'h30343667) * $signed(16'h0);
  assign twiddle4_1_235_imag = T20550 + T20548;
  assign T20548 = $signed(T20549) / $signed(22'h100000);
  assign T20549 = $signed(31'h2a3f5039) * $signed(16'hffff);
  assign T20550 = $signed(T20551) / $signed(22'h100000);
  assign T20551 = $signed(31'h301316ea) * $signed(16'h0);
  assign T20552 = T18725[1'h0:1'h0];
  assign T20553 = T18725[1'h1:1'h1];
  assign T20554 = T20575 ? T20565 : T20555;
  assign T20555 = T20564 ? twiddle4_1_237_imag : twiddle4_1_236_imag;
  assign twiddle4_1_236_imag = T20558 + T20556;
  assign T20556 = $signed(T20557) / $signed(22'h100000);
  assign T20557 = $signed(31'h2a650525) * $signed(16'hffff);
  assign T20558 = $signed(T20559) / $signed(22'h100000);
  assign T20559 = $signed(31'h2ff1d9c6) * $signed(16'h0);
  assign twiddle4_1_237_imag = T20562 + T20560;
  assign T20560 = $signed(T20561) / $signed(22'h100000);
  assign T20561 = $signed(31'h2a8a9fea) * $signed(16'hffff);
  assign T20562 = $signed(T20563) / $signed(22'h100000);
  assign T20563 = $signed(31'h2fd07f0f) * $signed(16'h0);
  assign T20564 = T18725[1'h0:1'h0];
  assign T20565 = T20574 ? twiddle4_1_239_imag : twiddle4_1_238_imag;
  assign twiddle4_1_238_imag = T20568 + T20566;
  assign T20566 = $signed(T20567) / $signed(22'h100000);
  assign T20567 = $signed(31'h2ab02071) * $signed(16'hffff);
  assign T20568 = $signed(T20569) / $signed(22'h100000);
  assign T20569 = $signed(31'h2faf06d9) * $signed(16'h0);
  assign twiddle4_1_239_imag = T20572 + T20570;
  assign T20570 = $signed(T20571) / $signed(22'h100000);
  assign T20571 = $signed(31'h2ad586a3) * $signed(16'hffff);
  assign T20572 = $signed(T20573) / $signed(22'h100000);
  assign T20573 = $signed(31'h2f8d7139) * $signed(16'h0);
  assign T20574 = T18725[1'h0:1'h0];
  assign T20575 = T18725[1'h1:1'h1];
  assign T20576 = T18725[2'h2:2'h2];
  assign T20577 = T18725[2'h3:2'h3];
  assign T20578 = T20671 ? T20625 : T20579;
  assign T20579 = T20624 ? T20602 : T20580;
  assign T20580 = T20601 ? T20591 : T20581;
  assign T20581 = T20590 ? twiddle4_1_241_imag : twiddle4_1_240_imag;
  assign twiddle4_1_240_imag = T20584 + T20582;
  assign T20582 = $signed(T20583) / $signed(22'h100000);
  assign T20583 = $signed(31'h2afad269) * $signed(16'hffff);
  assign T20584 = $signed(T20585) / $signed(22'h100000);
  assign T20585 = $signed(31'h2f6bbe44) * $signed(16'h0);
  assign twiddle4_1_241_imag = T20588 + T20586;
  assign T20586 = $signed(T20587) / $signed(22'h100000);
  assign T20587 = $signed(31'h2b2003ab) * $signed(16'hffff);
  assign T20588 = $signed(T20589) / $signed(22'h100000);
  assign T20589 = $signed(31'h2f49ee0f) * $signed(16'h0);
  assign T20590 = T18725[1'h0:1'h0];
  assign T20591 = T20600 ? twiddle4_1_243_imag : twiddle4_1_242_imag;
  assign twiddle4_1_242_imag = T20594 + T20592;
  assign T20592 = $signed(T20593) / $signed(22'h100000);
  assign T20593 = $signed(31'h2b451a54) * $signed(16'hffff);
  assign T20594 = $signed(T20595) / $signed(22'h100000);
  assign T20595 = $signed(31'h2f2800ae) * $signed(16'h0);
  assign twiddle4_1_243_imag = T20598 + T20596;
  assign T20596 = $signed(T20597) / $signed(22'h100000);
  assign T20597 = $signed(31'h2b6a164c) * $signed(16'hffff);
  assign T20598 = $signed(T20599) / $signed(22'h100000);
  assign T20599 = $signed(31'h2f05f637) * $signed(16'h0);
  assign T20600 = T18725[1'h0:1'h0];
  assign T20601 = T18725[1'h1:1'h1];
  assign T20602 = T20623 ? T20613 : T20603;
  assign T20603 = T20612 ? twiddle4_1_245_imag : twiddle4_1_244_imag;
  assign twiddle4_1_244_imag = T20606 + T20604;
  assign T20604 = $signed(T20605) / $signed(22'h100000);
  assign T20605 = $signed(31'h2b8ef77c) * $signed(16'hffff);
  assign T20606 = $signed(T20607) / $signed(22'h100000);
  assign T20607 = $signed(31'h2ee3cebe) * $signed(16'h0);
  assign twiddle4_1_245_imag = T20610 + T20608;
  assign T20608 = $signed(T20609) / $signed(22'h100000);
  assign T20609 = $signed(31'h2bb3bdce) * $signed(16'hffff);
  assign T20610 = $signed(T20611) / $signed(22'h100000);
  assign T20611 = $signed(31'h2ec18a58) * $signed(16'h0);
  assign T20612 = T18725[1'h0:1'h0];
  assign T20613 = T20622 ? twiddle4_1_247_imag : twiddle4_1_246_imag;
  assign twiddle4_1_246_imag = T20616 + T20614;
  assign T20614 = $signed(T20615) / $signed(22'h100000);
  assign T20615 = $signed(31'h2bd8692b) * $signed(16'hffff);
  assign T20616 = $signed(T20617) / $signed(22'h100000);
  assign T20617 = $signed(31'h2e9f291b) * $signed(16'h0);
  assign twiddle4_1_247_imag = T20620 + T20618;
  assign T20618 = $signed(T20619) / $signed(22'h100000);
  assign T20619 = $signed(31'h2bfcf97b) * $signed(16'hffff);
  assign T20620 = $signed(T20621) / $signed(22'h100000);
  assign T20621 = $signed(31'h2e7cab1c) * $signed(16'h0);
  assign T20622 = T18725[1'h0:1'h0];
  assign T20623 = T18725[1'h1:1'h1];
  assign T20624 = T18725[2'h2:2'h2];
  assign T20625 = T20670 ? T20648 : T20626;
  assign T20626 = T20647 ? T20637 : T20627;
  assign T20627 = T20636 ? twiddle4_1_249_imag : twiddle4_1_248_imag;
  assign twiddle4_1_248_imag = T20630 + T20628;
  assign T20628 = $signed(T20629) / $signed(22'h100000);
  assign T20629 = $signed(31'h2c216eaa) * $signed(16'hffff);
  assign T20630 = $signed(T20631) / $signed(22'h100000);
  assign T20631 = $signed(31'h2e5a106f) * $signed(16'h0);
  assign twiddle4_1_249_imag = T20634 + T20632;
  assign T20632 = $signed(T20633) / $signed(22'h100000);
  assign T20633 = $signed(31'h2c45c89f) * $signed(16'hffff);
  assign T20634 = $signed(T20635) / $signed(22'h100000);
  assign T20635 = $signed(31'h2e37592c) * $signed(16'h0);
  assign T20636 = T18725[1'h0:1'h0];
  assign T20637 = T20646 ? twiddle4_1_251_imag : twiddle4_1_250_imag;
  assign twiddle4_1_250_imag = T20640 + T20638;
  assign T20638 = $signed(T20639) / $signed(22'h100000);
  assign T20639 = $signed(31'h2c6a0746) * $signed(16'hffff);
  assign T20640 = $signed(T20641) / $signed(22'h100000);
  assign T20641 = $signed(31'h2e148566) * $signed(16'h0);
  assign twiddle4_1_251_imag = T20644 + T20642;
  assign T20642 = $signed(T20643) / $signed(22'h100000);
  assign T20643 = $signed(31'h2c8e2a86) * $signed(16'hffff);
  assign T20644 = $signed(T20645) / $signed(22'h100000);
  assign T20645 = $signed(31'h2df19533) * $signed(16'h0);
  assign T20646 = T18725[1'h0:1'h0];
  assign T20647 = T18725[1'h1:1'h1];
  assign T20648 = T20669 ? T20659 : T20649;
  assign T20649 = T20658 ? twiddle4_1_253_imag : twiddle4_1_252_imag;
  assign twiddle4_1_252_imag = T20652 + T20650;
  assign T20650 = $signed(T20651) / $signed(22'h100000);
  assign T20651 = $signed(31'h2cb2324b) * $signed(16'hffff);
  assign T20652 = $signed(T20653) / $signed(22'h100000);
  assign T20653 = $signed(31'h2dce88a9) * $signed(16'h0);
  assign twiddle4_1_253_imag = T20656 + T20654;
  assign T20654 = $signed(T20655) / $signed(22'h100000);
  assign T20655 = $signed(31'h2cd61e7e) * $signed(16'hffff);
  assign T20656 = $signed(T20657) / $signed(22'h100000);
  assign T20657 = $signed(31'h2dab5fde) * $signed(16'h0);
  assign T20658 = T18725[1'h0:1'h0];
  assign T20659 = T20668 ? twiddle4_1_255_imag : twiddle4_1_254_imag;
  assign twiddle4_1_254_imag = T20662 + T20660;
  assign T20660 = $signed(T20661) / $signed(22'h100000);
  assign T20661 = $signed(31'h2cf9ef09) * $signed(16'hffff);
  assign T20662 = $signed(T20663) / $signed(22'h100000);
  assign T20663 = $signed(31'h2d881ae7) * $signed(16'h0);
  assign twiddle4_1_255_imag = T20666 + T20664;
  assign T20664 = $signed(T20665) / $signed(22'h100000);
  assign T20665 = $signed(31'h2d1da3d5) * $signed(16'hffff);
  assign T20666 = $signed(T20667) / $signed(22'h100000);
  assign T20667 = $signed(31'h2d64b9da) * $signed(16'h0);
  assign T20668 = T18725[1'h0:1'h0];
  assign T20669 = T18725[1'h1:1'h1];
  assign T20670 = T18725[2'h2:2'h2];
  assign T20671 = T18725[2'h3:2'h3];
  assign T20672 = T18725[3'h4:3'h4];
  assign T20673 = T18725[3'h5:3'h5];
  assign T20674 = T18725[3'h6:3'h6];
  assign T20675 = T19823[6'h2e:6'h2e];
  assign T20676 = T18725[3'h7:3'h7];
  assign T20677 = {T22634, T20678};
  assign T20678 = T22633 ? T21529 : T20679;
  assign T20679 = T21528 ? T21062 : T20680;
  assign T20680 = T21061 ? T20871 : T20681;
  assign T20681 = T20870 ? T20776 : T20682;
  assign T20682 = T20775 ? T20729 : T20683;
  assign T20683 = T20728 ? T20706 : T20684;
  assign T20684 = T20705 ? T20695 : T20685;
  assign T20685 = T20694 ? twiddle4_1_257_imag : twiddle4_1_256_imag;
  assign twiddle4_1_256_imag = T20688 + T20686;
  assign T20686 = $signed(T20687) / $signed(22'h100000);
  assign T20687 = $signed(31'h2d413ccc) * $signed(16'hffff);
  assign T20688 = $signed(T20689) / $signed(22'h100000);
  assign T20689 = $signed(31'h2d413ccc) * $signed(16'h0);
  assign twiddle4_1_257_imag = T20692 + T20690;
  assign T20690 = $signed(T20691) / $signed(22'h100000);
  assign T20691 = $signed(31'h2d64b9da) * $signed(16'hffff);
  assign T20692 = $signed(T20693) / $signed(22'h100000);
  assign T20693 = $signed(31'h2d1da3d5) * $signed(16'h0);
  assign T20694 = T18725[1'h0:1'h0];
  assign T20695 = T20704 ? twiddle4_1_259_imag : twiddle4_1_258_imag;
  assign twiddle4_1_258_imag = T20698 + T20696;
  assign T20696 = $signed(T20697) / $signed(22'h100000);
  assign T20697 = $signed(31'h2d881ae7) * $signed(16'hffff);
  assign T20698 = $signed(T20699) / $signed(22'h100000);
  assign T20699 = $signed(31'h2cf9ef09) * $signed(16'h0);
  assign twiddle4_1_259_imag = T20702 + T20700;
  assign T20700 = $signed(T20701) / $signed(22'h100000);
  assign T20701 = $signed(31'h2dab5fde) * $signed(16'hffff);
  assign T20702 = $signed(T20703) / $signed(22'h100000);
  assign T20703 = $signed(31'h2cd61e7e) * $signed(16'h0);
  assign T20704 = T18725[1'h0:1'h0];
  assign T20705 = T18725[1'h1:1'h1];
  assign T20706 = T20727 ? T20717 : T20707;
  assign T20707 = T20716 ? twiddle4_1_261_imag : twiddle4_1_260_imag;
  assign twiddle4_1_260_imag = T20710 + T20708;
  assign T20708 = $signed(T20709) / $signed(22'h100000);
  assign T20709 = $signed(31'h2dce88a9) * $signed(16'hffff);
  assign T20710 = $signed(T20711) / $signed(22'h100000);
  assign T20711 = $signed(31'h2cb2324b) * $signed(16'h0);
  assign twiddle4_1_261_imag = T20714 + T20712;
  assign T20712 = $signed(T20713) / $signed(22'h100000);
  assign T20713 = $signed(31'h2df19533) * $signed(16'hffff);
  assign T20714 = $signed(T20715) / $signed(22'h100000);
  assign T20715 = $signed(31'h2c8e2a86) * $signed(16'h0);
  assign T20716 = T18725[1'h0:1'h0];
  assign T20717 = T20726 ? twiddle4_1_263_imag : twiddle4_1_262_imag;
  assign twiddle4_1_262_imag = T20720 + T20718;
  assign T20718 = $signed(T20719) / $signed(22'h100000);
  assign T20719 = $signed(31'h2e148566) * $signed(16'hffff);
  assign T20720 = $signed(T20721) / $signed(22'h100000);
  assign T20721 = $signed(31'h2c6a0746) * $signed(16'h0);
  assign twiddle4_1_263_imag = T20724 + T20722;
  assign T20722 = $signed(T20723) / $signed(22'h100000);
  assign T20723 = $signed(31'h2e37592c) * $signed(16'hffff);
  assign T20724 = $signed(T20725) / $signed(22'h100000);
  assign T20725 = $signed(31'h2c45c89f) * $signed(16'h0);
  assign T20726 = T18725[1'h0:1'h0];
  assign T20727 = T18725[1'h1:1'h1];
  assign T20728 = T18725[2'h2:2'h2];
  assign T20729 = T20774 ? T20752 : T20730;
  assign T20730 = T20751 ? T20741 : T20731;
  assign T20731 = T20740 ? twiddle4_1_265_imag : twiddle4_1_264_imag;
  assign twiddle4_1_264_imag = T20734 + T20732;
  assign T20732 = $signed(T20733) / $signed(22'h100000);
  assign T20733 = $signed(31'h2e5a106f) * $signed(16'hffff);
  assign T20734 = $signed(T20735) / $signed(22'h100000);
  assign T20735 = $signed(31'h2c216eaa) * $signed(16'h0);
  assign twiddle4_1_265_imag = T20738 + T20736;
  assign T20736 = $signed(T20737) / $signed(22'h100000);
  assign T20737 = $signed(31'h2e7cab1c) * $signed(16'hffff);
  assign T20738 = $signed(T20739) / $signed(22'h100000);
  assign T20739 = $signed(31'h2bfcf97b) * $signed(16'h0);
  assign T20740 = T18725[1'h0:1'h0];
  assign T20741 = T20750 ? twiddle4_1_267_imag : twiddle4_1_266_imag;
  assign twiddle4_1_266_imag = T20744 + T20742;
  assign T20742 = $signed(T20743) / $signed(22'h100000);
  assign T20743 = $signed(31'h2e9f291b) * $signed(16'hffff);
  assign T20744 = $signed(T20745) / $signed(22'h100000);
  assign T20745 = $signed(31'h2bd8692b) * $signed(16'h0);
  assign twiddle4_1_267_imag = T20748 + T20746;
  assign T20746 = $signed(T20747) / $signed(22'h100000);
  assign T20747 = $signed(31'h2ec18a58) * $signed(16'hffff);
  assign T20748 = $signed(T20749) / $signed(22'h100000);
  assign T20749 = $signed(31'h2bb3bdce) * $signed(16'h0);
  assign T20750 = T18725[1'h0:1'h0];
  assign T20751 = T18725[1'h1:1'h1];
  assign T20752 = T20773 ? T20763 : T20753;
  assign T20753 = T20762 ? twiddle4_1_269_imag : twiddle4_1_268_imag;
  assign twiddle4_1_268_imag = T20756 + T20754;
  assign T20754 = $signed(T20755) / $signed(22'h100000);
  assign T20755 = $signed(31'h2ee3cebe) * $signed(16'hffff);
  assign T20756 = $signed(T20757) / $signed(22'h100000);
  assign T20757 = $signed(31'h2b8ef77c) * $signed(16'h0);
  assign twiddle4_1_269_imag = T20760 + T20758;
  assign T20758 = $signed(T20759) / $signed(22'h100000);
  assign T20759 = $signed(31'h2f05f637) * $signed(16'hffff);
  assign T20760 = $signed(T20761) / $signed(22'h100000);
  assign T20761 = $signed(31'h2b6a164c) * $signed(16'h0);
  assign T20762 = T18725[1'h0:1'h0];
  assign T20763 = T20772 ? twiddle4_1_271_imag : twiddle4_1_270_imag;
  assign twiddle4_1_270_imag = T20766 + T20764;
  assign T20764 = $signed(T20765) / $signed(22'h100000);
  assign T20765 = $signed(31'h2f2800ae) * $signed(16'hffff);
  assign T20766 = $signed(T20767) / $signed(22'h100000);
  assign T20767 = $signed(31'h2b451a54) * $signed(16'h0);
  assign twiddle4_1_271_imag = T20770 + T20768;
  assign T20768 = $signed(T20769) / $signed(22'h100000);
  assign T20769 = $signed(31'h2f49ee0f) * $signed(16'hffff);
  assign T20770 = $signed(T20771) / $signed(22'h100000);
  assign T20771 = $signed(31'h2b2003ab) * $signed(16'h0);
  assign T20772 = T18725[1'h0:1'h0];
  assign T20773 = T18725[1'h1:1'h1];
  assign T20774 = T18725[2'h2:2'h2];
  assign T20775 = T18725[2'h3:2'h3];
  assign T20776 = T20869 ? T20823 : T20777;
  assign T20777 = T20822 ? T20800 : T20778;
  assign T20778 = T20799 ? T20789 : T20779;
  assign T20779 = T20788 ? twiddle4_1_273_imag : twiddle4_1_272_imag;
  assign twiddle4_1_272_imag = T20782 + T20780;
  assign T20780 = $signed(T20781) / $signed(22'h100000);
  assign T20781 = $signed(31'h2f6bbe44) * $signed(16'hffff);
  assign T20782 = $signed(T20783) / $signed(22'h100000);
  assign T20783 = $signed(31'h2afad269) * $signed(16'h0);
  assign twiddle4_1_273_imag = T20786 + T20784;
  assign T20784 = $signed(T20785) / $signed(22'h100000);
  assign T20785 = $signed(31'h2f8d7139) * $signed(16'hffff);
  assign T20786 = $signed(T20787) / $signed(22'h100000);
  assign T20787 = $signed(31'h2ad586a3) * $signed(16'h0);
  assign T20788 = T18725[1'h0:1'h0];
  assign T20789 = T20798 ? twiddle4_1_275_imag : twiddle4_1_274_imag;
  assign twiddle4_1_274_imag = T20792 + T20790;
  assign T20790 = $signed(T20791) / $signed(22'h100000);
  assign T20791 = $signed(31'h2faf06d9) * $signed(16'hffff);
  assign T20792 = $signed(T20793) / $signed(22'h100000);
  assign T20793 = $signed(31'h2ab02071) * $signed(16'h0);
  assign twiddle4_1_275_imag = T20796 + T20794;
  assign T20794 = $signed(T20795) / $signed(22'h100000);
  assign T20795 = $signed(31'h2fd07f0f) * $signed(16'hffff);
  assign T20796 = $signed(T20797) / $signed(22'h100000);
  assign T20797 = $signed(31'h2a8a9fea) * $signed(16'h0);
  assign T20798 = T18725[1'h0:1'h0];
  assign T20799 = T18725[1'h1:1'h1];
  assign T20800 = T20821 ? T20811 : T20801;
  assign T20801 = T20810 ? twiddle4_1_277_imag : twiddle4_1_276_imag;
  assign twiddle4_1_276_imag = T20804 + T20802;
  assign T20802 = $signed(T20803) / $signed(22'h100000);
  assign T20803 = $signed(31'h2ff1d9c6) * $signed(16'hffff);
  assign T20804 = $signed(T20805) / $signed(22'h100000);
  assign T20805 = $signed(31'h2a650525) * $signed(16'h0);
  assign twiddle4_1_277_imag = T20808 + T20806;
  assign T20806 = $signed(T20807) / $signed(22'h100000);
  assign T20807 = $signed(31'h301316ea) * $signed(16'hffff);
  assign T20808 = $signed(T20809) / $signed(22'h100000);
  assign T20809 = $signed(31'h2a3f5039) * $signed(16'h0);
  assign T20810 = T18725[1'h0:1'h0];
  assign T20811 = T20820 ? twiddle4_1_279_imag : twiddle4_1_278_imag;
  assign twiddle4_1_278_imag = T20814 + T20812;
  assign T20812 = $signed(T20813) / $signed(22'h100000);
  assign T20813 = $signed(31'h30343667) * $signed(16'hffff);
  assign T20814 = $signed(T20815) / $signed(22'h100000);
  assign T20815 = $signed(31'h2a19813e) * $signed(16'h0);
  assign twiddle4_1_279_imag = T20818 + T20816;
  assign T20816 = $signed(T20817) / $signed(22'h100000);
  assign T20817 = $signed(31'h30553827) * $signed(16'hffff);
  assign T20818 = $signed(T20819) / $signed(22'h100000);
  assign T20819 = $signed(31'h29f3984b) * $signed(16'h0);
  assign T20820 = T18725[1'h0:1'h0];
  assign T20821 = T18725[1'h1:1'h1];
  assign T20822 = T18725[2'h2:2'h2];
  assign T20823 = T20868 ? T20846 : T20824;
  assign T20824 = T20845 ? T20835 : T20825;
  assign T20825 = T20834 ? twiddle4_1_281_imag : twiddle4_1_280_imag;
  assign twiddle4_1_280_imag = T20828 + T20826;
  assign T20826 = $signed(T20827) / $signed(22'h100000);
  assign T20827 = $signed(31'h30761c17) * $signed(16'hffff);
  assign T20828 = $signed(T20829) / $signed(22'h100000);
  assign T20829 = $signed(31'h29cd9577) * $signed(16'h0);
  assign twiddle4_1_281_imag = T20832 + T20830;
  assign T20830 = $signed(T20831) / $signed(22'h100000);
  assign T20831 = $signed(31'h3096e223) * $signed(16'hffff);
  assign T20832 = $signed(T20833) / $signed(22'h100000);
  assign T20833 = $signed(31'h29a778da) * $signed(16'h0);
  assign T20834 = T18725[1'h0:1'h0];
  assign T20835 = T20844 ? twiddle4_1_283_imag : twiddle4_1_282_imag;
  assign twiddle4_1_282_imag = T20838 + T20836;
  assign T20836 = $signed(T20837) / $signed(22'h100000);
  assign T20837 = $signed(31'h30b78a35) * $signed(16'hffff);
  assign T20838 = $signed(T20839) / $signed(22'h100000);
  assign T20839 = $signed(31'h2981428b) * $signed(16'h0);
  assign twiddle4_1_283_imag = T20842 + T20840;
  assign T20840 = $signed(T20841) / $signed(22'h100000);
  assign T20841 = $signed(31'h30d8143b) * $signed(16'hffff);
  assign T20842 = $signed(T20843) / $signed(22'h100000);
  assign T20843 = $signed(31'h295af2a2) * $signed(16'h0);
  assign T20844 = T18725[1'h0:1'h0];
  assign T20845 = T18725[1'h1:1'h1];
  assign T20846 = T20867 ? T20857 : T20847;
  assign T20847 = T20856 ? twiddle4_1_285_imag : twiddle4_1_284_imag;
  assign twiddle4_1_284_imag = T20850 + T20848;
  assign T20848 = $signed(T20849) / $signed(22'h100000);
  assign T20849 = $signed(31'h30f8801f) * $signed(16'hffff);
  assign T20850 = $signed(T20851) / $signed(22'h100000);
  assign T20851 = $signed(31'h29348937) * $signed(16'h0);
  assign twiddle4_1_285_imag = T20854 + T20852;
  assign T20852 = $signed(T20853) / $signed(22'h100000);
  assign T20853 = $signed(31'h3118cdce) * $signed(16'hffff);
  assign T20854 = $signed(T20855) / $signed(22'h100000);
  assign T20855 = $signed(31'h290e0660) * $signed(16'h0);
  assign T20856 = T18725[1'h0:1'h0];
  assign T20857 = T20866 ? twiddle4_1_287_imag : twiddle4_1_286_imag;
  assign twiddle4_1_286_imag = T20860 + T20858;
  assign T20858 = $signed(T20859) / $signed(22'h100000);
  assign T20859 = $signed(31'h3138fd34) * $signed(16'hffff);
  assign T20860 = $signed(T20861) / $signed(22'h100000);
  assign T20861 = $signed(31'h28e76a37) * $signed(16'h0);
  assign twiddle4_1_287_imag = T20864 + T20862;
  assign T20862 = $signed(T20863) / $signed(22'h100000);
  assign T20863 = $signed(31'h31590e3d) * $signed(16'hffff);
  assign T20864 = $signed(T20865) / $signed(22'h100000);
  assign T20865 = $signed(31'h28c0b4d2) * $signed(16'h0);
  assign T20866 = T18725[1'h0:1'h0];
  assign T20867 = T18725[1'h1:1'h1];
  assign T20868 = T18725[2'h2:2'h2];
  assign T20869 = T18725[2'h3:2'h3];
  assign T20870 = T18725[3'h4:3'h4];
  assign T20871 = T21060 ? T20966 : T20872;
  assign T20872 = T20965 ? T20919 : T20873;
  assign T20873 = T20918 ? T20896 : T20874;
  assign T20874 = T20895 ? T20885 : T20875;
  assign T20875 = T20884 ? twiddle4_1_289_imag : twiddle4_1_288_imag;
  assign twiddle4_1_288_imag = T20878 + T20876;
  assign T20876 = $signed(T20877) / $signed(22'h100000);
  assign T20877 = $signed(31'h317900d6) * $signed(16'hffff);
  assign T20878 = $signed(T20879) / $signed(22'h100000);
  assign T20879 = $signed(31'h2899e64a) * $signed(16'h0);
  assign twiddle4_1_289_imag = T20882 + T20880;
  assign T20880 = $signed(T20881) / $signed(22'h100000);
  assign T20881 = $signed(31'h3198d4ea) * $signed(16'hffff);
  assign T20882 = $signed(T20883) / $signed(22'h100000);
  assign T20883 = $signed(31'h2872feb6) * $signed(16'h0);
  assign T20884 = T18725[1'h0:1'h0];
  assign T20885 = T20894 ? twiddle4_1_291_imag : twiddle4_1_290_imag;
  assign twiddle4_1_290_imag = T20888 + T20886;
  assign T20886 = $signed(T20887) / $signed(22'h100000);
  assign T20887 = $signed(31'h31b88a66) * $signed(16'hffff);
  assign T20888 = $signed(T20889) / $signed(22'h100000);
  assign T20889 = $signed(31'h284bfe2f) * $signed(16'h0);
  assign twiddle4_1_291_imag = T20892 + T20890;
  assign T20890 = $signed(T20891) / $signed(22'h100000);
  assign T20891 = $signed(31'h31d82136) * $signed(16'hffff);
  assign T20892 = $signed(T20893) / $signed(22'h100000);
  assign T20893 = $signed(31'h2824e4cc) * $signed(16'h0);
  assign T20894 = T18725[1'h0:1'h0];
  assign T20895 = T18725[1'h1:1'h1];
  assign T20896 = T20917 ? T20907 : T20897;
  assign T20897 = T20906 ? twiddle4_1_293_imag : twiddle4_1_292_imag;
  assign twiddle4_1_292_imag = T20900 + T20898;
  assign T20898 = $signed(T20899) / $signed(22'h100000);
  assign T20899 = $signed(31'h31f79947) * $signed(16'hffff);
  assign T20900 = $signed(T20901) / $signed(22'h100000);
  assign T20901 = $signed(31'h27fdb2a6) * $signed(16'h0);
  assign twiddle4_1_293_imag = T20904 + T20902;
  assign T20902 = $signed(T20903) / $signed(22'h100000);
  assign T20903 = $signed(31'h3216f286) * $signed(16'hffff);
  assign T20904 = $signed(T20905) / $signed(22'h100000);
  assign T20905 = $signed(31'h27d667d5) * $signed(16'h0);
  assign T20906 = T18725[1'h0:1'h0];
  assign T20907 = T20916 ? twiddle4_1_295_imag : twiddle4_1_294_imag;
  assign twiddle4_1_294_imag = T20910 + T20908;
  assign T20908 = $signed(T20909) / $signed(22'h100000);
  assign T20909 = $signed(31'h32362cdf) * $signed(16'hffff);
  assign T20910 = $signed(T20911) / $signed(22'h100000);
  assign T20911 = $signed(31'h27af0471) * $signed(16'h0);
  assign twiddle4_1_295_imag = T20914 + T20912;
  assign T20912 = $signed(T20913) / $signed(22'h100000);
  assign T20913 = $signed(31'h3255483f) * $signed(16'hffff);
  assign T20914 = $signed(T20915) / $signed(22'h100000);
  assign T20915 = $signed(31'h27878893) * $signed(16'h0);
  assign T20916 = T18725[1'h0:1'h0];
  assign T20917 = T18725[1'h1:1'h1];
  assign T20918 = T18725[2'h2:2'h2];
  assign T20919 = T20964 ? T20942 : T20920;
  assign T20920 = T20941 ? T20931 : T20921;
  assign T20921 = T20930 ? twiddle4_1_297_imag : twiddle4_1_296_imag;
  assign twiddle4_1_296_imag = T20924 + T20922;
  assign T20922 = $signed(T20923) / $signed(22'h100000);
  assign T20923 = $signed(31'h32744493) * $signed(16'hffff);
  assign T20924 = $signed(T20925) / $signed(22'h100000);
  assign T20925 = $signed(31'h275ff452) * $signed(16'h0);
  assign twiddle4_1_297_imag = T20928 + T20926;
  assign T20926 = $signed(T20927) / $signed(22'h100000);
  assign T20927 = $signed(31'h329321c7) * $signed(16'hffff);
  assign T20928 = $signed(T20929) / $signed(22'h100000);
  assign T20929 = $signed(31'h273847c7) * $signed(16'h0);
  assign T20930 = T18725[1'h0:1'h0];
  assign T20931 = T20940 ? twiddle4_1_299_imag : twiddle4_1_298_imag;
  assign twiddle4_1_298_imag = T20934 + T20932;
  assign T20932 = $signed(T20933) / $signed(22'h100000);
  assign T20933 = $signed(31'h32b1dfc9) * $signed(16'hffff);
  assign T20934 = $signed(T20935) / $signed(22'h100000);
  assign T20935 = $signed(31'h2710830b) * $signed(16'h0);
  assign twiddle4_1_299_imag = T20938 + T20936;
  assign T20936 = $signed(T20937) / $signed(22'h100000);
  assign T20937 = $signed(31'h32d07e85) * $signed(16'hffff);
  assign T20938 = $signed(T20939) / $signed(22'h100000);
  assign T20939 = $signed(31'h26e8a637) * $signed(16'h0);
  assign T20940 = T18725[1'h0:1'h0];
  assign T20941 = T18725[1'h1:1'h1];
  assign T20942 = T20963 ? T20953 : T20943;
  assign T20943 = T20952 ? twiddle4_1_301_imag : twiddle4_1_300_imag;
  assign twiddle4_1_300_imag = T20946 + T20944;
  assign T20944 = $signed(T20945) / $signed(22'h100000);
  assign T20945 = $signed(31'h32eefde9) * $signed(16'hffff);
  assign T20946 = $signed(T20947) / $signed(22'h100000);
  assign T20947 = $signed(31'h26c0b162) * $signed(16'h0);
  assign twiddle4_1_301_imag = T20950 + T20948;
  assign T20948 = $signed(T20949) / $signed(22'h100000);
  assign T20949 = $signed(31'h330d5de2) * $signed(16'hffff);
  assign T20950 = $signed(T20951) / $signed(22'h100000);
  assign T20951 = $signed(31'h2698a4a5) * $signed(16'h0);
  assign T20952 = T18725[1'h0:1'h0];
  assign T20953 = T20962 ? twiddle4_1_303_imag : twiddle4_1_302_imag;
  assign twiddle4_1_302_imag = T20956 + T20954;
  assign T20954 = $signed(T20955) / $signed(22'h100000);
  assign T20955 = $signed(31'h332b9e5d) * $signed(16'hffff);
  assign T20956 = $signed(T20957) / $signed(22'h100000);
  assign T20957 = $signed(31'h2670801a) * $signed(16'h0);
  assign twiddle4_1_303_imag = T20960 + T20958;
  assign T20958 = $signed(T20959) / $signed(22'h100000);
  assign T20959 = $signed(31'h3349bf48) * $signed(16'hffff);
  assign T20960 = $signed(T20961) / $signed(22'h100000);
  assign T20961 = $signed(31'h264843d8) * $signed(16'h0);
  assign T20962 = T18725[1'h0:1'h0];
  assign T20963 = T18725[1'h1:1'h1];
  assign T20964 = T18725[2'h2:2'h2];
  assign T20965 = T18725[2'h3:2'h3];
  assign T20966 = T21059 ? T21013 : T20967;
  assign T20967 = T21012 ? T20990 : T20968;
  assign T20968 = T20989 ? T20979 : T20969;
  assign T20969 = T20978 ? twiddle4_1_305_imag : twiddle4_1_304_imag;
  assign twiddle4_1_304_imag = T20972 + T20970;
  assign T20970 = $signed(T20971) / $signed(22'h100000);
  assign T20971 = $signed(31'h3367c08f) * $signed(16'hffff);
  assign T20972 = $signed(T20973) / $signed(22'h100000);
  assign T20973 = $signed(31'h261feff9) * $signed(16'h0);
  assign twiddle4_1_305_imag = T20976 + T20974;
  assign T20974 = $signed(T20975) / $signed(22'h100000);
  assign T20975 = $signed(31'h3385a221) * $signed(16'hffff);
  assign T20976 = $signed(T20977) / $signed(22'h100000);
  assign T20977 = $signed(31'h25f78496) * $signed(16'h0);
  assign T20978 = T18725[1'h0:1'h0];
  assign T20979 = T20988 ? twiddle4_1_307_imag : twiddle4_1_306_imag;
  assign twiddle4_1_306_imag = T20982 + T20980;
  assign T20980 = $signed(T20981) / $signed(22'h100000);
  assign T20981 = $signed(31'h33a363eb) * $signed(16'hffff);
  assign T20982 = $signed(T20983) / $signed(22'h100000);
  assign T20983 = $signed(31'h25cf01c7) * $signed(16'h0);
  assign twiddle4_1_307_imag = T20986 + T20984;
  assign T20984 = $signed(T20985) / $signed(22'h100000);
  assign T20985 = $signed(31'h33c105db) * $signed(16'hffff);
  assign T20986 = $signed(T20987) / $signed(22'h100000);
  assign T20987 = $signed(31'h25a667a6) * $signed(16'h0);
  assign T20988 = T18725[1'h0:1'h0];
  assign T20989 = T18725[1'h1:1'h1];
  assign T20990 = T21011 ? T21001 : T20991;
  assign T20991 = T21000 ? twiddle4_1_309_imag : twiddle4_1_308_imag;
  assign twiddle4_1_308_imag = T20994 + T20992;
  assign T20992 = $signed(T20993) / $signed(22'h100000);
  assign T20993 = $signed(31'h33de87de) * $signed(16'hffff);
  assign T20994 = $signed(T20995) / $signed(22'h100000);
  assign T20995 = $signed(31'h257db64b) * $signed(16'h0);
  assign twiddle4_1_309_imag = T20998 + T20996;
  assign T20996 = $signed(T20997) / $signed(22'h100000);
  assign T20997 = $signed(31'h33fbe9e2) * $signed(16'hffff);
  assign T20998 = $signed(T20999) / $signed(22'h100000);
  assign T20999 = $signed(31'h2554edd0) * $signed(16'h0);
  assign T21000 = T18725[1'h0:1'h0];
  assign T21001 = T21010 ? twiddle4_1_311_imag : twiddle4_1_310_imag;
  assign twiddle4_1_310_imag = T21004 + T21002;
  assign T21002 = $signed(T21003) / $signed(22'h100000);
  assign T21003 = $signed(31'h34192bd5) * $signed(16'hffff);
  assign T21004 = $signed(T21005) / $signed(22'h100000);
  assign T21005 = $signed(31'h252c0e4e) * $signed(16'h0);
  assign twiddle4_1_311_imag = T21008 + T21006;
  assign T21006 = $signed(T21007) / $signed(22'h100000);
  assign T21007 = $signed(31'h34364da5) * $signed(16'hffff);
  assign T21008 = $signed(T21009) / $signed(22'h100000);
  assign T21009 = $signed(31'h250317de) * $signed(16'h0);
  assign T21010 = T18725[1'h0:1'h0];
  assign T21011 = T18725[1'h1:1'h1];
  assign T21012 = T18725[2'h2:2'h2];
  assign T21013 = T21058 ? T21036 : T21014;
  assign T21014 = T21035 ? T21025 : T21015;
  assign T21015 = T21024 ? twiddle4_1_313_imag : twiddle4_1_312_imag;
  assign twiddle4_1_312_imag = T21018 + T21016;
  assign T21016 = $signed(T21017) / $signed(22'h100000);
  assign T21017 = $signed(31'h34534f40) * $signed(16'hffff);
  assign T21018 = $signed(T21019) / $signed(22'h100000);
  assign T21019 = $signed(31'h24da0a99) * $signed(16'h0);
  assign twiddle4_1_313_imag = T21022 + T21020;
  assign T21020 = $signed(T21021) / $signed(22'h100000);
  assign T21021 = $signed(31'h34703094) * $signed(16'hffff);
  assign T21022 = $signed(T21023) / $signed(22'h100000);
  assign T21023 = $signed(31'h24b0e699) * $signed(16'h0);
  assign T21024 = T18725[1'h0:1'h0];
  assign T21025 = T21034 ? twiddle4_1_315_imag : twiddle4_1_314_imag;
  assign twiddle4_1_314_imag = T21028 + T21026;
  assign T21026 = $signed(T21027) / $signed(22'h100000);
  assign T21027 = $signed(31'h348cf190) * $signed(16'hffff);
  assign T21028 = $signed(T21029) / $signed(22'h100000);
  assign T21029 = $signed(31'h2487abf7) * $signed(16'h0);
  assign twiddle4_1_315_imag = T21032 + T21030;
  assign T21030 = $signed(T21031) / $signed(22'h100000);
  assign T21031 = $signed(31'h34a99221) * $signed(16'hffff);
  assign T21032 = $signed(T21033) / $signed(22'h100000);
  assign T21033 = $signed(31'h245e5acc) * $signed(16'h0);
  assign T21034 = T18725[1'h0:1'h0];
  assign T21035 = T18725[1'h1:1'h1];
  assign T21036 = T21057 ? T21047 : T21037;
  assign T21037 = T21046 ? twiddle4_1_317_imag : twiddle4_1_316_imag;
  assign twiddle4_1_316_imag = T21040 + T21038;
  assign T21038 = $signed(T21039) / $signed(22'h100000);
  assign T21039 = $signed(31'h34c61236) * $signed(16'hffff);
  assign T21040 = $signed(T21041) / $signed(22'h100000);
  assign T21041 = $signed(31'h2434f332) * $signed(16'h0);
  assign twiddle4_1_317_imag = T21044 + T21042;
  assign T21042 = $signed(T21043) / $signed(22'h100000);
  assign T21043 = $signed(31'h34e271bd) * $signed(16'hffff);
  assign T21044 = $signed(T21045) / $signed(22'h100000);
  assign T21045 = $signed(31'h240b7542) * $signed(16'h0);
  assign T21046 = T18725[1'h0:1'h0];
  assign T21047 = T21056 ? twiddle4_1_319_imag : twiddle4_1_318_imag;
  assign twiddle4_1_318_imag = T21050 + T21048;
  assign T21048 = $signed(T21049) / $signed(22'h100000);
  assign T21049 = $signed(31'h34feb0a5) * $signed(16'hffff);
  assign T21050 = $signed(T21051) / $signed(22'h100000);
  assign T21051 = $signed(31'h23e1e117) * $signed(16'h0);
  assign twiddle4_1_319_imag = T21054 + T21052;
  assign T21052 = $signed(T21053) / $signed(22'h100000);
  assign T21053 = $signed(31'h351acedc) * $signed(16'hffff);
  assign T21054 = $signed(T21055) / $signed(22'h100000);
  assign T21055 = $signed(31'h23b836c9) * $signed(16'h0);
  assign T21056 = T18725[1'h0:1'h0];
  assign T21057 = T18725[1'h1:1'h1];
  assign T21058 = T18725[2'h2:2'h2];
  assign T21059 = T18725[2'h3:2'h3];
  assign T21060 = T18725[3'h4:3'h4];
  assign T21061 = T18725[3'h5:3'h5];
  assign T21062 = T21527 ? T21273 : T21063;
  assign T21063 = T21272 ? T21158 : T21064;
  assign T21064 = T21157 ? T21111 : T21065;
  assign T21065 = T21110 ? T21088 : T21066;
  assign T21066 = T21087 ? T21077 : T21067;
  assign T21067 = T21076 ? twiddle4_1_321_imag : twiddle4_1_320_imag;
  assign twiddle4_1_320_imag = T21070 + T21068;
  assign T21068 = $signed(T21069) / $signed(22'h100000);
  assign T21069 = $signed(31'h3536cc52) * $signed(16'hffff);
  assign T21070 = $signed(T21071) / $signed(22'h100000);
  assign T21071 = $signed(31'h238e7673) * $signed(16'h0);
  assign twiddle4_1_321_imag = T21074 + T21072;
  assign T21072 = $signed(T21073) / $signed(22'h100000);
  assign T21073 = $signed(31'h3552a8f4) * $signed(16'hffff);
  assign T21074 = $signed(T21075) / $signed(22'h100000);
  assign T21075 = $signed(31'h2364a02e) * $signed(16'h0);
  assign T21076 = T18725[1'h0:1'h0];
  assign T21077 = T21086 ? twiddle4_1_323_imag : twiddle4_1_322_imag;
  assign twiddle4_1_322_imag = T21080 + T21078;
  assign T21078 = $signed(T21079) / $signed(22'h100000);
  assign T21079 = $signed(31'h356e64b2) * $signed(16'hffff);
  assign T21080 = $signed(T21081) / $signed(22'h100000);
  assign T21081 = $signed(31'h233ab413) * $signed(16'h0);
  assign twiddle4_1_323_imag = T21084 + T21082;
  assign T21082 = $signed(T21083) / $signed(22'h100000);
  assign T21083 = $signed(31'h3589ff7a) * $signed(16'hffff);
  assign T21084 = $signed(T21085) / $signed(22'h100000);
  assign T21085 = $signed(31'h2310b23e) * $signed(16'h0);
  assign T21086 = T18725[1'h0:1'h0];
  assign T21087 = T18725[1'h1:1'h1];
  assign T21088 = T21109 ? T21099 : T21089;
  assign T21089 = T21098 ? twiddle4_1_325_imag : twiddle4_1_324_imag;
  assign twiddle4_1_324_imag = T21092 + T21090;
  assign T21090 = $signed(T21091) / $signed(22'h100000);
  assign T21091 = $signed(31'h35a5793c) * $signed(16'hffff);
  assign T21092 = $signed(T21093) / $signed(22'h100000);
  assign T21093 = $signed(31'h22e69ac7) * $signed(16'h0);
  assign twiddle4_1_325_imag = T21096 + T21094;
  assign T21094 = $signed(T21095) / $signed(22'h100000);
  assign T21095 = $signed(31'h35c0d1e6) * $signed(16'hffff);
  assign T21096 = $signed(T21097) / $signed(22'h100000);
  assign T21097 = $signed(31'h22bc6dc9) * $signed(16'h0);
  assign T21098 = T18725[1'h0:1'h0];
  assign T21099 = T21108 ? twiddle4_1_327_imag : twiddle4_1_326_imag;
  assign twiddle4_1_326_imag = T21102 + T21100;
  assign T21100 = $signed(T21101) / $signed(22'h100000);
  assign T21101 = $signed(31'h35dc0968) * $signed(16'hffff);
  assign T21102 = $signed(T21103) / $signed(22'h100000);
  assign T21103 = $signed(31'h22922b5e) * $signed(16'h0);
  assign twiddle4_1_327_imag = T21106 + T21104;
  assign T21104 = $signed(T21105) / $signed(22'h100000);
  assign T21105 = $signed(31'h35f71fb1) * $signed(16'hffff);
  assign T21106 = $signed(T21107) / $signed(22'h100000);
  assign T21107 = $signed(31'h2267d39f) * $signed(16'h0);
  assign T21108 = T18725[1'h0:1'h0];
  assign T21109 = T18725[1'h1:1'h1];
  assign T21110 = T18725[2'h2:2'h2];
  assign T21111 = T21156 ? T21134 : T21112;
  assign T21112 = T21133 ? T21123 : T21113;
  assign T21113 = T21122 ? twiddle4_1_329_imag : twiddle4_1_328_imag;
  assign twiddle4_1_328_imag = T21116 + T21114;
  assign T21114 = $signed(T21115) / $signed(22'h100000);
  assign T21115 = $signed(31'h361214b0) * $signed(16'hffff);
  assign T21116 = $signed(T21117) / $signed(22'h100000);
  assign T21117 = $signed(31'h223d66a8) * $signed(16'h0);
  assign twiddle4_1_329_imag = T21120 + T21118;
  assign T21118 = $signed(T21119) / $signed(22'h100000);
  assign T21119 = $signed(31'h362ce854) * $signed(16'hffff);
  assign T21120 = $signed(T21121) / $signed(22'h100000);
  assign T21121 = $signed(31'h2212e491) * $signed(16'h0);
  assign T21122 = T18725[1'h0:1'h0];
  assign T21123 = T21132 ? twiddle4_1_331_imag : twiddle4_1_330_imag;
  assign twiddle4_1_330_imag = T21126 + T21124;
  assign T21124 = $signed(T21125) / $signed(22'h100000);
  assign T21125 = $signed(31'h36479a8e) * $signed(16'hffff);
  assign T21126 = $signed(T21127) / $signed(22'h100000);
  assign T21127 = $signed(31'h21e84d76) * $signed(16'h0);
  assign twiddle4_1_331_imag = T21130 + T21128;
  assign T21128 = $signed(T21129) / $signed(22'h100000);
  assign T21129 = $signed(31'h36622b4b) * $signed(16'hffff);
  assign T21130 = $signed(T21131) / $signed(22'h100000);
  assign T21131 = $signed(31'h21bda170) * $signed(16'h0);
  assign T21132 = T18725[1'h0:1'h0];
  assign T21133 = T18725[1'h1:1'h1];
  assign T21134 = T21155 ? T21145 : T21135;
  assign T21135 = T21144 ? twiddle4_1_333_imag : twiddle4_1_332_imag;
  assign twiddle4_1_332_imag = T21138 + T21136;
  assign T21136 = $signed(T21137) / $signed(22'h100000);
  assign T21137 = $signed(31'h367c9a7d) * $signed(16'hffff);
  assign T21138 = $signed(T21139) / $signed(22'h100000);
  assign T21139 = $signed(31'h2192e09a) * $signed(16'h0);
  assign twiddle4_1_333_imag = T21142 + T21140;
  assign T21140 = $signed(T21141) / $signed(22'h100000);
  assign T21141 = $signed(31'h3696e813) * $signed(16'hffff);
  assign T21142 = $signed(T21143) / $signed(22'h100000);
  assign T21143 = $signed(31'h21680b0f) * $signed(16'h0);
  assign T21144 = T18725[1'h0:1'h0];
  assign T21145 = T21154 ? twiddle4_1_335_imag : twiddle4_1_334_imag;
  assign twiddle4_1_334_imag = T21148 + T21146;
  assign T21146 = $signed(T21147) / $signed(22'h100000);
  assign T21147 = $signed(31'h36b113fd) * $signed(16'hffff);
  assign T21148 = $signed(T21149) / $signed(22'h100000);
  assign T21149 = $signed(31'h213d20e8) * $signed(16'h0);
  assign twiddle4_1_335_imag = T21152 + T21150;
  assign T21150 = $signed(T21151) / $signed(22'h100000);
  assign T21151 = $signed(31'h36cb1e29) * $signed(16'hffff);
  assign T21152 = $signed(T21153) / $signed(22'h100000);
  assign T21153 = $signed(31'h21122240) * $signed(16'h0);
  assign T21154 = T18725[1'h0:1'h0];
  assign T21155 = T18725[1'h1:1'h1];
  assign T21156 = T18725[2'h2:2'h2];
  assign T21157 = T18725[2'h3:2'h3];
  assign T21158 = T21271 ? T21209 : T21159;
  assign T21159 = T21208 ? T21182 : T21160;
  assign T21160 = T21181 ? T21171 : T21161;
  assign T21161 = T21170 ? twiddle4_1_337_imag : twiddle4_1_336_imag;
  assign twiddle4_1_336_imag = T21164 + T21162;
  assign T21162 = $signed(T21163) / $signed(22'h100000);
  assign T21163 = $signed(31'h36e5068a) * $signed(16'hffff);
  assign T21164 = $signed(T21165) / $signed(22'h100000);
  assign T21165 = $signed(31'h20e70f32) * $signed(16'h0);
  assign twiddle4_1_337_imag = T21168 + T21166;
  assign T21166 = $signed(T21167) / $signed(22'h100000);
  assign T21167 = $signed(31'h36fecd0d) * $signed(16'hffff);
  assign T21168 = $signed(T21169) / $signed(22'h100000);
  assign T21169 = $signed(31'h20bbe7d8) * $signed(16'h0);
  assign T21170 = T18725[1'h0:1'h0];
  assign T21171 = T21180 ? twiddle4_1_339_imag : twiddle4_1_338_imag;
  assign twiddle4_1_338_imag = T21174 + T21172;
  assign T21172 = $signed(T21173) / $signed(22'h100000);
  assign T21173 = $signed(31'h371871a4) * $signed(16'hffff);
  assign T21174 = $signed(T21175) / $signed(22'h100000);
  assign T21175 = $signed(31'h2090ac4d) * $signed(16'h0);
  assign twiddle4_1_339_imag = T21178 + T21176;
  assign T21176 = $signed(T21177) / $signed(22'h100000);
  assign T21177 = $signed(31'h3731f43f) * $signed(16'hffff);
  assign T21178 = $signed(T21179) / $signed(22'h100000);
  assign T21179 = $signed(31'h20655cab) * $signed(16'h0);
  assign T21180 = T18725[1'h0:1'h0];
  assign T21181 = T18725[1'h1:1'h1];
  assign T21182 = T21207 ? T21193 : T21183;
  assign T21183 = T21192 ? twiddle4_1_341_imag : twiddle4_1_340_imag;
  assign twiddle4_1_340_imag = T21186 + T21184;
  assign T21184 = $signed(T21185) / $signed(22'h100000);
  assign T21185 = $signed(31'h374b54ce) * $signed(16'hffff);
  assign T21186 = $signed(T21187) / $signed(22'h100000);
  assign T21187 = $signed(31'h2039f90e) * $signed(16'h0);
  assign twiddle4_1_341_imag = T21190 + T21188;
  assign T21188 = $signed(T21189) / $signed(22'h100000);
  assign T21189 = $signed(31'h37649341) * $signed(16'hffff);
  assign T21190 = $signed(T21191) / $signed(22'h100000);
  assign T21191 = $signed(31'h200e8190) * $signed(16'h0);
  assign T21192 = T18725[1'h0:1'h0];
  assign T21193 = T21206 ? twiddle4_1_343_imag : twiddle4_1_342_imag;
  assign twiddle4_1_342_imag = T21196 + T21194;
  assign T21194 = $signed(T21195) / $signed(22'h100000);
  assign T21195 = $signed(31'h377daf89) * $signed(16'hffff);
  assign T21196 = {T21199, T21197};
  assign T21197 = $signed(T21198) / $signed(22'h100000);
  assign T21198 = $signed(30'h1fe2f64b) * $signed(16'h0);
  assign T21199 = T21197[6'h2d:6'h2d];
  assign twiddle4_1_343_imag = T21202 + T21200;
  assign T21200 = $signed(T21201) / $signed(22'h100000);
  assign T21201 = $signed(31'h3796a996) * $signed(16'hffff);
  assign T21202 = {T21205, T21203};
  assign T21203 = $signed(T21204) / $signed(22'h100000);
  assign T21204 = $signed(30'h1fb7575c) * $signed(16'h0);
  assign T21205 = T21203[6'h2d:6'h2d];
  assign T21206 = T18725[1'h0:1'h0];
  assign T21207 = T18725[1'h1:1'h1];
  assign T21208 = T18725[2'h2:2'h2];
  assign T21209 = T21270 ? T21240 : T21210;
  assign T21210 = T21239 ? T21225 : T21211;
  assign T21211 = T21224 ? twiddle4_1_345_imag : twiddle4_1_344_imag;
  assign twiddle4_1_344_imag = T21214 + T21212;
  assign T21212 = $signed(T21213) / $signed(22'h100000);
  assign T21213 = $signed(31'h37af8158) * $signed(16'hffff);
  assign T21214 = {T21217, T21215};
  assign T21215 = $signed(T21216) / $signed(22'h100000);
  assign T21216 = $signed(30'h1f8ba4db) * $signed(16'h0);
  assign T21217 = T21215[6'h2d:6'h2d];
  assign twiddle4_1_345_imag = T21220 + T21218;
  assign T21218 = $signed(T21219) / $signed(22'h100000);
  assign T21219 = $signed(31'h37c836c2) * $signed(16'hffff);
  assign T21220 = {T21223, T21221};
  assign T21221 = $signed(T21222) / $signed(22'h100000);
  assign T21222 = $signed(30'h1f5fdee6) * $signed(16'h0);
  assign T21223 = T21221[6'h2d:6'h2d];
  assign T21224 = T18725[1'h0:1'h0];
  assign T21225 = T21238 ? twiddle4_1_347_imag : twiddle4_1_346_imag;
  assign twiddle4_1_346_imag = T21228 + T21226;
  assign T21226 = $signed(T21227) / $signed(22'h100000);
  assign T21227 = $signed(31'h37e0c9c2) * $signed(16'hffff);
  assign T21228 = {T21231, T21229};
  assign T21229 = $signed(T21230) / $signed(22'h100000);
  assign T21230 = $signed(30'h1f340596) * $signed(16'h0);
  assign T21231 = T21229[6'h2d:6'h2d];
  assign twiddle4_1_347_imag = T21234 + T21232;
  assign T21232 = $signed(T21233) / $signed(22'h100000);
  assign T21233 = $signed(31'h37f93a4b) * $signed(16'hffff);
  assign T21234 = {T21237, T21235};
  assign T21235 = $signed(T21236) / $signed(22'h100000);
  assign T21236 = $signed(30'h1f081906) * $signed(16'h0);
  assign T21237 = T21235[6'h2d:6'h2d];
  assign T21238 = T18725[1'h0:1'h0];
  assign T21239 = T18725[1'h1:1'h1];
  assign T21240 = T21269 ? T21255 : T21241;
  assign T21241 = T21254 ? twiddle4_1_349_imag : twiddle4_1_348_imag;
  assign twiddle4_1_348_imag = T21244 + T21242;
  assign T21242 = $signed(T21243) / $signed(22'h100000);
  assign T21243 = $signed(31'h3811884c) * $signed(16'hffff);
  assign T21244 = {T21247, T21245};
  assign T21245 = $signed(T21246) / $signed(22'h100000);
  assign T21246 = $signed(30'h1edc1952) * $signed(16'h0);
  assign T21247 = T21245[6'h2d:6'h2d];
  assign twiddle4_1_349_imag = T21250 + T21248;
  assign T21248 = $signed(T21249) / $signed(22'h100000);
  assign T21249 = $signed(31'h3829b3b8) * $signed(16'hffff);
  assign T21250 = {T21253, T21251};
  assign T21251 = $signed(T21252) / $signed(22'h100000);
  assign T21252 = $signed(30'h1eb00695) * $signed(16'h0);
  assign T21253 = T21251[6'h2d:6'h2d];
  assign T21254 = T18725[1'h0:1'h0];
  assign T21255 = T21268 ? twiddle4_1_351_imag : twiddle4_1_350_imag;
  assign twiddle4_1_350_imag = T21258 + T21256;
  assign T21256 = $signed(T21257) / $signed(22'h100000);
  assign T21257 = $signed(31'h3841bc7f) * $signed(16'hffff);
  assign T21258 = {T21261, T21259};
  assign T21259 = $signed(T21260) / $signed(22'h100000);
  assign T21260 = $signed(30'h1e83e0ea) * $signed(16'h0);
  assign T21261 = T21259[6'h2d:6'h2d];
  assign twiddle4_1_351_imag = T21264 + T21262;
  assign T21262 = $signed(T21263) / $signed(22'h100000);
  assign T21263 = $signed(31'h3859a292) * $signed(16'hffff);
  assign T21264 = {T21267, T21265};
  assign T21265 = $signed(T21266) / $signed(22'h100000);
  assign T21266 = $signed(30'h1e57a86d) * $signed(16'h0);
  assign T21267 = T21265[6'h2d:6'h2d];
  assign T21268 = T18725[1'h0:1'h0];
  assign T21269 = T18725[1'h1:1'h1];
  assign T21270 = T18725[2'h2:2'h2];
  assign T21271 = T18725[2'h3:2'h3];
  assign T21272 = T18725[3'h4:3'h4];
  assign T21273 = T21526 ? T21400 : T21274;
  assign T21274 = T21399 ? T21337 : T21275;
  assign T21275 = T21336 ? T21306 : T21276;
  assign T21276 = T21305 ? T21291 : T21277;
  assign T21277 = T21290 ? twiddle4_1_353_imag : twiddle4_1_352_imag;
  assign twiddle4_1_352_imag = T21280 + T21278;
  assign T21278 = $signed(T21279) / $signed(22'h100000);
  assign T21279 = $signed(31'h387165e3) * $signed(16'hffff);
  assign T21280 = {T21283, T21281};
  assign T21281 = $signed(T21282) / $signed(22'h100000);
  assign T21282 = $signed(30'h1e2b5d38) * $signed(16'h0);
  assign T21283 = T21281[6'h2d:6'h2d];
  assign twiddle4_1_353_imag = T21286 + T21284;
  assign T21284 = $signed(T21285) / $signed(22'h100000);
  assign T21285 = $signed(31'h38890662) * $signed(16'hffff);
  assign T21286 = {T21289, T21287};
  assign T21287 = $signed(T21288) / $signed(22'h100000);
  assign T21288 = $signed(30'h1dfeff66) * $signed(16'h0);
  assign T21289 = T21287[6'h2d:6'h2d];
  assign T21290 = T18725[1'h0:1'h0];
  assign T21291 = T21304 ? twiddle4_1_355_imag : twiddle4_1_354_imag;
  assign twiddle4_1_354_imag = T21294 + T21292;
  assign T21292 = $signed(T21293) / $signed(22'h100000);
  assign T21293 = $signed(31'h38a08402) * $signed(16'hffff);
  assign T21294 = {T21297, T21295};
  assign T21295 = $signed(T21296) / $signed(22'h100000);
  assign T21296 = $signed(30'h1dd28f14) * $signed(16'h0);
  assign T21297 = T21295[6'h2d:6'h2d];
  assign twiddle4_1_355_imag = T21300 + T21298;
  assign T21298 = $signed(T21299) / $signed(22'h100000);
  assign T21299 = $signed(31'h38b7deb3) * $signed(16'hffff);
  assign T21300 = {T21303, T21301};
  assign T21301 = $signed(T21302) / $signed(22'h100000);
  assign T21302 = $signed(30'h1da60c5c) * $signed(16'h0);
  assign T21303 = T21301[6'h2d:6'h2d];
  assign T21304 = T18725[1'h0:1'h0];
  assign T21305 = T18725[1'h1:1'h1];
  assign T21306 = T21335 ? T21321 : T21307;
  assign T21307 = T21320 ? twiddle4_1_357_imag : twiddle4_1_356_imag;
  assign twiddle4_1_356_imag = T21310 + T21308;
  assign T21308 = $signed(T21309) / $signed(22'h100000);
  assign T21309 = $signed(31'h38cf1669) * $signed(16'hffff);
  assign T21310 = {T21313, T21311};
  assign T21311 = $signed(T21312) / $signed(22'h100000);
  assign T21312 = $signed(30'h1d79775b) * $signed(16'h0);
  assign T21313 = T21311[6'h2d:6'h2d];
  assign twiddle4_1_357_imag = T21316 + T21314;
  assign T21314 = $signed(T21315) / $signed(22'h100000);
  assign T21315 = $signed(31'h38e62b13) * $signed(16'hffff);
  assign T21316 = {T21319, T21317};
  assign T21317 = $signed(T21318) / $signed(22'h100000);
  assign T21318 = $signed(30'h1d4cd02b) * $signed(16'h0);
  assign T21319 = T21317[6'h2d:6'h2d];
  assign T21320 = T18725[1'h0:1'h0];
  assign T21321 = T21334 ? twiddle4_1_359_imag : twiddle4_1_358_imag;
  assign twiddle4_1_358_imag = T21324 + T21322;
  assign T21322 = $signed(T21323) / $signed(22'h100000);
  assign T21323 = $signed(31'h38fd1ca4) * $signed(16'hffff);
  assign T21324 = {T21327, T21325};
  assign T21325 = $signed(T21326) / $signed(22'h100000);
  assign T21326 = $signed(30'h1d2016e8) * $signed(16'h0);
  assign T21327 = T21325[6'h2d:6'h2d];
  assign twiddle4_1_359_imag = T21330 + T21328;
  assign T21328 = $signed(T21329) / $signed(22'h100000);
  assign T21329 = $signed(31'h3913eb0e) * $signed(16'hffff);
  assign T21330 = {T21333, T21331};
  assign T21331 = $signed(T21332) / $signed(22'h100000);
  assign T21332 = $signed(30'h1cf34bae) * $signed(16'h0);
  assign T21333 = T21331[6'h2d:6'h2d];
  assign T21334 = T18725[1'h0:1'h0];
  assign T21335 = T18725[1'h1:1'h1];
  assign T21336 = T18725[2'h2:2'h2];
  assign T21337 = T21398 ? T21368 : T21338;
  assign T21338 = T21367 ? T21353 : T21339;
  assign T21339 = T21352 ? twiddle4_1_361_imag : twiddle4_1_360_imag;
  assign twiddle4_1_360_imag = T21342 + T21340;
  assign T21340 = $signed(T21341) / $signed(22'h100000);
  assign T21341 = $signed(31'h392a9642) * $signed(16'hffff);
  assign T21342 = {T21345, T21343};
  assign T21343 = $signed(T21344) / $signed(22'h100000);
  assign T21344 = $signed(30'h1cc66e99) * $signed(16'h0);
  assign T21345 = T21343[6'h2d:6'h2d];
  assign twiddle4_1_361_imag = T21348 + T21346;
  assign T21346 = $signed(T21347) / $signed(22'h100000);
  assign T21347 = $signed(31'h39411e33) * $signed(16'hffff);
  assign T21348 = {T21351, T21349};
  assign T21349 = $signed(T21350) / $signed(22'h100000);
  assign T21350 = $signed(30'h1c997fc3) * $signed(16'h0);
  assign T21351 = T21349[6'h2d:6'h2d];
  assign T21352 = T18725[1'h0:1'h0];
  assign T21353 = T21366 ? twiddle4_1_363_imag : twiddle4_1_362_imag;
  assign twiddle4_1_362_imag = T21356 + T21354;
  assign T21354 = $signed(T21355) / $signed(22'h100000);
  assign T21355 = $signed(31'h395782d3) * $signed(16'hffff);
  assign T21356 = {T21359, T21357};
  assign T21357 = $signed(T21358) / $signed(22'h100000);
  assign T21358 = $signed(30'h1c6c7f49) * $signed(16'h0);
  assign T21359 = T21357[6'h2d:6'h2d];
  assign twiddle4_1_363_imag = T21362 + T21360;
  assign T21360 = $signed(T21361) / $signed(22'h100000);
  assign T21361 = $signed(31'h396dc414) * $signed(16'hffff);
  assign T21362 = {T21365, T21363};
  assign T21363 = $signed(T21364) / $signed(22'h100000);
  assign T21364 = $signed(30'h1c3f6d47) * $signed(16'h0);
  assign T21365 = T21363[6'h2d:6'h2d];
  assign T21366 = T18725[1'h0:1'h0];
  assign T21367 = T18725[1'h1:1'h1];
  assign T21368 = T21397 ? T21383 : T21369;
  assign T21369 = T21382 ? twiddle4_1_365_imag : twiddle4_1_364_imag;
  assign twiddle4_1_364_imag = T21372 + T21370;
  assign T21370 = $signed(T21371) / $signed(22'h100000);
  assign T21371 = $signed(31'h3983e1e7) * $signed(16'hffff);
  assign T21372 = {T21375, T21373};
  assign T21373 = $signed(T21374) / $signed(22'h100000);
  assign T21374 = $signed(30'h1c1249d8) * $signed(16'h0);
  assign T21375 = T21373[6'h2d:6'h2d];
  assign twiddle4_1_365_imag = T21378 + T21376;
  assign T21376 = $signed(T21377) / $signed(22'h100000);
  assign T21377 = $signed(31'h3999dc41) * $signed(16'hffff);
  assign T21378 = {T21381, T21379};
  assign T21379 = $signed(T21380) / $signed(22'h100000);
  assign T21380 = $signed(30'h1be51517) * $signed(16'h0);
  assign T21381 = T21379[6'h2d:6'h2d];
  assign T21382 = T18725[1'h0:1'h0];
  assign T21383 = T21396 ? twiddle4_1_367_imag : twiddle4_1_366_imag;
  assign twiddle4_1_366_imag = T21386 + T21384;
  assign T21384 = $signed(T21385) / $signed(22'h100000);
  assign T21385 = $signed(31'h39afb313) * $signed(16'hffff);
  assign T21386 = {T21389, T21387};
  assign T21387 = $signed(T21388) / $signed(22'h100000);
  assign T21388 = $signed(30'h1bb7cf23) * $signed(16'h0);
  assign T21389 = T21387[6'h2d:6'h2d];
  assign twiddle4_1_367_imag = T21392 + T21390;
  assign T21390 = $signed(T21391) / $signed(22'h100000);
  assign T21391 = $signed(31'h39c5664f) * $signed(16'hffff);
  assign T21392 = {T21395, T21393};
  assign T21393 = $signed(T21394) / $signed(22'h100000);
  assign T21394 = $signed(30'h1b8a7814) * $signed(16'h0);
  assign T21395 = T21393[6'h2d:6'h2d];
  assign T21396 = T18725[1'h0:1'h0];
  assign T21397 = T18725[1'h1:1'h1];
  assign T21398 = T18725[2'h2:2'h2];
  assign T21399 = T18725[2'h3:2'h3];
  assign T21400 = T21525 ? T21463 : T21401;
  assign T21401 = T21462 ? T21432 : T21402;
  assign T21402 = T21431 ? T21417 : T21403;
  assign T21403 = T21416 ? twiddle4_1_369_imag : twiddle4_1_368_imag;
  assign twiddle4_1_368_imag = T21406 + T21404;
  assign T21404 = $signed(T21405) / $signed(22'h100000);
  assign T21405 = $signed(31'h39daf5e8) * $signed(16'hffff);
  assign T21406 = {T21409, T21407};
  assign T21407 = $signed(T21408) / $signed(22'h100000);
  assign T21408 = $signed(30'h1b5d1009) * $signed(16'h0);
  assign T21409 = T21407[6'h2d:6'h2d];
  assign twiddle4_1_369_imag = T21412 + T21410;
  assign T21410 = $signed(T21411) / $signed(22'h100000);
  assign T21411 = $signed(31'h39f061d1) * $signed(16'hffff);
  assign T21412 = {T21415, T21413};
  assign T21413 = $signed(T21414) / $signed(22'h100000);
  assign T21414 = $signed(30'h1b2f971d) * $signed(16'h0);
  assign T21415 = T21413[6'h2d:6'h2d];
  assign T21416 = T18725[1'h0:1'h0];
  assign T21417 = T21430 ? twiddle4_1_371_imag : twiddle4_1_370_imag;
  assign twiddle4_1_370_imag = T21420 + T21418;
  assign T21418 = $signed(T21419) / $signed(22'h100000);
  assign T21419 = $signed(31'h3a05a9fd) * $signed(16'hffff);
  assign T21420 = {T21423, T21421};
  assign T21421 = $signed(T21422) / $signed(22'h100000);
  assign T21422 = $signed(30'h1b020d6c) * $signed(16'h0);
  assign T21423 = T21421[6'h2d:6'h2d];
  assign twiddle4_1_371_imag = T21426 + T21424;
  assign T21424 = $signed(T21425) / $signed(22'h100000);
  assign T21425 = $signed(31'h3a1ace5e) * $signed(16'hffff);
  assign T21426 = {T21429, T21427};
  assign T21427 = $signed(T21428) / $signed(22'h100000);
  assign T21428 = $signed(30'h1ad47312) * $signed(16'h0);
  assign T21429 = T21427[6'h2d:6'h2d];
  assign T21430 = T18725[1'h0:1'h0];
  assign T21431 = T18725[1'h1:1'h1];
  assign T21432 = T21461 ? T21447 : T21433;
  assign T21433 = T21446 ? twiddle4_1_373_imag : twiddle4_1_372_imag;
  assign twiddle4_1_372_imag = T21436 + T21434;
  assign T21434 = $signed(T21435) / $signed(22'h100000);
  assign T21435 = $signed(31'h3a2fcee8) * $signed(16'hffff);
  assign T21436 = {T21439, T21437};
  assign T21437 = $signed(T21438) / $signed(22'h100000);
  assign T21438 = $signed(30'h1aa6c82b) * $signed(16'h0);
  assign T21439 = T21437[6'h2d:6'h2d];
  assign twiddle4_1_373_imag = T21442 + T21440;
  assign T21440 = $signed(T21441) / $signed(22'h100000);
  assign T21441 = $signed(31'h3a44ab8d) * $signed(16'hffff);
  assign T21442 = {T21445, T21443};
  assign T21443 = $signed(T21444) / $signed(22'h100000);
  assign T21444 = $signed(30'h1a790cd3) * $signed(16'h0);
  assign T21445 = T21443[6'h2d:6'h2d];
  assign T21446 = T18725[1'h0:1'h0];
  assign T21447 = T21460 ? twiddle4_1_375_imag : twiddle4_1_374_imag;
  assign twiddle4_1_374_imag = T21450 + T21448;
  assign T21448 = $signed(T21449) / $signed(22'h100000);
  assign T21449 = $signed(31'h3a596441) * $signed(16'hffff);
  assign T21450 = {T21453, T21451};
  assign T21451 = $signed(T21452) / $signed(22'h100000);
  assign T21452 = $signed(30'h1a4b4127) * $signed(16'h0);
  assign T21453 = T21451[6'h2d:6'h2d];
  assign twiddle4_1_375_imag = T21456 + T21454;
  assign T21454 = $signed(T21455) / $signed(22'h100000);
  assign T21455 = $signed(31'h3a6df8f7) * $signed(16'hffff);
  assign T21456 = {T21459, T21457};
  assign T21457 = $signed(T21458) / $signed(22'h100000);
  assign T21458 = $signed(30'h1a1d6543) * $signed(16'h0);
  assign T21459 = T21457[6'h2d:6'h2d];
  assign T21460 = T18725[1'h0:1'h0];
  assign T21461 = T18725[1'h1:1'h1];
  assign T21462 = T18725[2'h2:2'h2];
  assign T21463 = T21524 ? T21494 : T21464;
  assign T21464 = T21493 ? T21479 : T21465;
  assign T21465 = T21478 ? twiddle4_1_377_imag : twiddle4_1_376_imag;
  assign twiddle4_1_376_imag = T21468 + T21466;
  assign T21466 = $signed(T21467) / $signed(22'h100000);
  assign T21467 = $signed(31'h3a8269a2) * $signed(16'hffff);
  assign T21468 = {T21471, T21469};
  assign T21469 = $signed(T21470) / $signed(22'h100000);
  assign T21470 = $signed(30'h19ef7943) * $signed(16'h0);
  assign T21471 = T21469[6'h2d:6'h2d];
  assign twiddle4_1_377_imag = T21474 + T21472;
  assign T21472 = $signed(T21473) / $signed(22'h100000);
  assign T21473 = $signed(31'h3a96b636) * $signed(16'hffff);
  assign T21474 = {T21477, T21475};
  assign T21475 = $signed(T21476) / $signed(22'h100000);
  assign T21476 = $signed(30'h19c17d44) * $signed(16'h0);
  assign T21477 = T21475[6'h2d:6'h2d];
  assign T21478 = T18725[1'h0:1'h0];
  assign T21479 = T21492 ? twiddle4_1_379_imag : twiddle4_1_378_imag;
  assign twiddle4_1_378_imag = T21482 + T21480;
  assign T21480 = $signed(T21481) / $signed(22'h100000);
  assign T21481 = $signed(31'h3aaadea5) * $signed(16'hffff);
  assign T21482 = {T21485, T21483};
  assign T21483 = $signed(T21484) / $signed(22'h100000);
  assign T21484 = $signed(30'h19937161) * $signed(16'h0);
  assign T21485 = T21483[6'h2d:6'h2d];
  assign twiddle4_1_379_imag = T21488 + T21486;
  assign T21486 = $signed(T21487) / $signed(22'h100000);
  assign T21487 = $signed(31'h3abee2e5) * $signed(16'hffff);
  assign T21488 = {T21491, T21489};
  assign T21489 = $signed(T21490) / $signed(22'h100000);
  assign T21490 = $signed(30'h196555b7) * $signed(16'h0);
  assign T21491 = T21489[6'h2d:6'h2d];
  assign T21492 = T18725[1'h0:1'h0];
  assign T21493 = T18725[1'h1:1'h1];
  assign T21494 = T21523 ? T21509 : T21495;
  assign T21495 = T21508 ? twiddle4_1_381_imag : twiddle4_1_380_imag;
  assign twiddle4_1_380_imag = T21498 + T21496;
  assign T21496 = $signed(T21497) / $signed(22'h100000);
  assign T21497 = $signed(31'h3ad2c2e7) * $signed(16'hffff);
  assign T21498 = {T21501, T21499};
  assign T21499 = $signed(T21500) / $signed(22'h100000);
  assign T21500 = $signed(30'h19372a63) * $signed(16'h0);
  assign T21501 = T21499[6'h2d:6'h2d];
  assign twiddle4_1_381_imag = T21504 + T21502;
  assign T21502 = $signed(T21503) / $signed(22'h100000);
  assign T21503 = $signed(31'h3ae67ea1) * $signed(16'hffff);
  assign T21504 = {T21507, T21505};
  assign T21505 = $signed(T21506) / $signed(22'h100000);
  assign T21506 = $signed(30'h1908ef81) * $signed(16'h0);
  assign T21507 = T21505[6'h2d:6'h2d];
  assign T21508 = T18725[1'h0:1'h0];
  assign T21509 = T21522 ? twiddle4_1_383_imag : twiddle4_1_382_imag;
  assign twiddle4_1_382_imag = T21512 + T21510;
  assign T21510 = $signed(T21511) / $signed(22'h100000);
  assign T21511 = $signed(31'h3afa1605) * $signed(16'hffff);
  assign T21512 = {T21515, T21513};
  assign T21513 = $signed(T21514) / $signed(22'h100000);
  assign T21514 = $signed(30'h18daa52e) * $signed(16'h0);
  assign T21515 = T21513[6'h2d:6'h2d];
  assign twiddle4_1_383_imag = T21518 + T21516;
  assign T21516 = $signed(T21517) / $signed(22'h100000);
  assign T21517 = $signed(31'h3b0d8908) * $signed(16'hffff);
  assign T21518 = {T21521, T21519};
  assign T21519 = $signed(T21520) / $signed(22'h100000);
  assign T21520 = $signed(30'h18ac4b86) * $signed(16'h0);
  assign T21521 = T21519[6'h2d:6'h2d];
  assign T21522 = T18725[1'h0:1'h0];
  assign T21523 = T18725[1'h1:1'h1];
  assign T21524 = T18725[2'h2:2'h2];
  assign T21525 = T18725[2'h3:2'h3];
  assign T21526 = T18725[3'h4:3'h4];
  assign T21527 = T18725[3'h5:3'h5];
  assign T21528 = T18725[3'h6:3'h6];
  assign T21529 = T22632 ? T22058 : T21530;
  assign T21530 = T22057 ? T21785 : T21531;
  assign T21531 = T21784 ? T21658 : T21532;
  assign T21532 = T21657 ? T21595 : T21533;
  assign T21533 = T21594 ? T21564 : T21534;
  assign T21534 = T21563 ? T21549 : T21535;
  assign T21535 = T21548 ? twiddle4_1_385_imag : twiddle4_1_384_imag;
  assign twiddle4_1_384_imag = T21538 + T21536;
  assign T21536 = $signed(T21537) / $signed(22'h100000);
  assign T21537 = $signed(31'h3b20d79e) * $signed(16'hffff);
  assign T21538 = {T21541, T21539};
  assign T21539 = $signed(T21540) / $signed(22'h100000);
  assign T21540 = $signed(30'h187de2a6) * $signed(16'h0);
  assign T21541 = T21539[6'h2d:6'h2d];
  assign twiddle4_1_385_imag = T21544 + T21542;
  assign T21542 = $signed(T21543) / $signed(22'h100000);
  assign T21543 = $signed(31'h3b3401bb) * $signed(16'hffff);
  assign T21544 = {T21547, T21545};
  assign T21545 = $signed(T21546) / $signed(22'h100000);
  assign T21546 = $signed(30'h184f6aaa) * $signed(16'h0);
  assign T21547 = T21545[6'h2d:6'h2d];
  assign T21548 = T18725[1'h0:1'h0];
  assign T21549 = T21562 ? twiddle4_1_387_imag : twiddle4_1_386_imag;
  assign twiddle4_1_386_imag = T21552 + T21550;
  assign T21550 = $signed(T21551) / $signed(22'h100000);
  assign T21551 = $signed(31'h3b470752) * $signed(16'hffff);
  assign T21552 = {T21555, T21553};
  assign T21553 = $signed(T21554) / $signed(22'h100000);
  assign T21554 = $signed(30'h1820e3b0) * $signed(16'h0);
  assign T21555 = T21553[6'h2d:6'h2d];
  assign twiddle4_1_387_imag = T21558 + T21556;
  assign T21556 = $signed(T21557) / $signed(22'h100000);
  assign T21557 = $signed(31'h3b59e859) * $signed(16'hffff);
  assign T21558 = {T21561, T21559};
  assign T21559 = $signed(T21560) / $signed(22'h100000);
  assign T21560 = $signed(30'h17f24dd3) * $signed(16'h0);
  assign T21561 = T21559[6'h2d:6'h2d];
  assign T21562 = T18725[1'h0:1'h0];
  assign T21563 = T18725[1'h1:1'h1];
  assign T21564 = T21593 ? T21579 : T21565;
  assign T21565 = T21578 ? twiddle4_1_389_imag : twiddle4_1_388_imag;
  assign twiddle4_1_388_imag = T21568 + T21566;
  assign T21566 = $signed(T21567) / $signed(22'h100000);
  assign T21567 = $signed(31'h3b6ca4c4) * $signed(16'hffff);
  assign T21568 = {T21571, T21569};
  assign T21569 = $signed(T21570) / $signed(22'h100000);
  assign T21570 = $signed(30'h17c3a931) * $signed(16'h0);
  assign T21571 = T21569[6'h2d:6'h2d];
  assign twiddle4_1_389_imag = T21574 + T21572;
  assign T21572 = $signed(T21573) / $signed(22'h100000);
  assign T21573 = $signed(31'h3b7f3c87) * $signed(16'hffff);
  assign T21574 = {T21577, T21575};
  assign T21575 = $signed(T21576) / $signed(22'h100000);
  assign T21576 = $signed(30'h1794f5e6) * $signed(16'h0);
  assign T21577 = T21575[6'h2d:6'h2d];
  assign T21578 = T18725[1'h0:1'h0];
  assign T21579 = T21592 ? twiddle4_1_391_imag : twiddle4_1_390_imag;
  assign twiddle4_1_390_imag = T21582 + T21580;
  assign T21580 = $signed(T21581) / $signed(22'h100000);
  assign T21581 = $signed(31'h3b91af96) * $signed(16'hffff);
  assign T21582 = {T21585, T21583};
  assign T21583 = $signed(T21584) / $signed(22'h100000);
  assign T21584 = $signed(30'h1766340f) * $signed(16'h0);
  assign T21585 = T21583[6'h2d:6'h2d];
  assign twiddle4_1_391_imag = T21588 + T21586;
  assign T21586 = $signed(T21587) / $signed(22'h100000);
  assign T21587 = $signed(31'h3ba3fde7) * $signed(16'hffff);
  assign T21588 = {T21591, T21589};
  assign T21589 = $signed(T21590) / $signed(22'h100000);
  assign T21590 = $signed(30'h173763c9) * $signed(16'h0);
  assign T21591 = T21589[6'h2d:6'h2d];
  assign T21592 = T18725[1'h0:1'h0];
  assign T21593 = T18725[1'h1:1'h1];
  assign T21594 = T18725[2'h2:2'h2];
  assign T21595 = T21656 ? T21626 : T21596;
  assign T21596 = T21625 ? T21611 : T21597;
  assign T21597 = T21610 ? twiddle4_1_393_imag : twiddle4_1_392_imag;
  assign twiddle4_1_392_imag = T21600 + T21598;
  assign T21598 = $signed(T21599) / $signed(22'h100000);
  assign T21599 = $signed(31'h3bb6276d) * $signed(16'hffff);
  assign T21600 = {T21603, T21601};
  assign T21601 = $signed(T21602) / $signed(22'h100000);
  assign T21602 = $signed(30'h17088530) * $signed(16'h0);
  assign T21603 = T21601[6'h2d:6'h2d];
  assign twiddle4_1_393_imag = T21606 + T21604;
  assign T21604 = $signed(T21605) / $signed(22'h100000);
  assign T21605 = $signed(31'h3bc82c1e) * $signed(16'hffff);
  assign T21606 = {T21609, T21607};
  assign T21607 = $signed(T21608) / $signed(22'h100000);
  assign T21608 = $signed(30'h16d99863) * $signed(16'h0);
  assign T21609 = T21607[6'h2d:6'h2d];
  assign T21610 = T18725[1'h0:1'h0];
  assign T21611 = T21624 ? twiddle4_1_395_imag : twiddle4_1_394_imag;
  assign twiddle4_1_394_imag = T21614 + T21612;
  assign T21612 = $signed(T21613) / $signed(22'h100000);
  assign T21613 = $signed(31'h3bda0bef) * $signed(16'hffff);
  assign T21614 = {T21617, T21615};
  assign T21615 = $signed(T21616) / $signed(22'h100000);
  assign T21616 = $signed(30'h16aa9d7d) * $signed(16'h0);
  assign T21617 = T21615[6'h2d:6'h2d];
  assign twiddle4_1_395_imag = T21620 + T21618;
  assign T21618 = $signed(T21619) / $signed(22'h100000);
  assign T21619 = $signed(31'h3bebc6d5) * $signed(16'hffff);
  assign T21620 = {T21623, T21621};
  assign T21621 = $signed(T21622) / $signed(22'h100000);
  assign T21622 = $signed(30'h167b949c) * $signed(16'h0);
  assign T21623 = T21621[6'h2d:6'h2d];
  assign T21624 = T18725[1'h0:1'h0];
  assign T21625 = T18725[1'h1:1'h1];
  assign T21626 = T21655 ? T21641 : T21627;
  assign T21627 = T21640 ? twiddle4_1_397_imag : twiddle4_1_396_imag;
  assign twiddle4_1_396_imag = T21630 + T21628;
  assign T21628 = $signed(T21629) / $signed(22'h100000);
  assign T21629 = $signed(31'h3bfd5cc4) * $signed(16'hffff);
  assign T21630 = {T21633, T21631};
  assign T21631 = $signed(T21632) / $signed(22'h100000);
  assign T21632 = $signed(30'h164c7ddd) * $signed(16'h0);
  assign T21633 = T21631[6'h2d:6'h2d];
  assign twiddle4_1_397_imag = T21636 + T21634;
  assign T21634 = $signed(T21635) / $signed(22'h100000);
  assign T21635 = $signed(31'h3c0ecdb2) * $signed(16'hffff);
  assign T21636 = {T21639, T21637};
  assign T21637 = $signed(T21638) / $signed(22'h100000);
  assign T21638 = $signed(30'h161d595c) * $signed(16'h0);
  assign T21639 = T21637[6'h2d:6'h2d];
  assign T21640 = T18725[1'h0:1'h0];
  assign T21641 = T21654 ? twiddle4_1_399_imag : twiddle4_1_398_imag;
  assign twiddle4_1_398_imag = T21644 + T21642;
  assign T21642 = $signed(T21643) / $signed(22'h100000);
  assign T21643 = $signed(31'h3c201994) * $signed(16'hffff);
  assign T21644 = {T21647, T21645};
  assign T21645 = $signed(T21646) / $signed(22'h100000);
  assign T21646 = $signed(30'h15ee2737) * $signed(16'h0);
  assign T21647 = T21645[6'h2d:6'h2d];
  assign twiddle4_1_399_imag = T21650 + T21648;
  assign T21648 = $signed(T21649) / $signed(22'h100000);
  assign T21649 = $signed(31'h3c31405f) * $signed(16'hffff);
  assign T21650 = {T21653, T21651};
  assign T21651 = $signed(T21652) / $signed(22'h100000);
  assign T21652 = $signed(30'h15bee78b) * $signed(16'h0);
  assign T21653 = T21651[6'h2d:6'h2d];
  assign T21654 = T18725[1'h0:1'h0];
  assign T21655 = T18725[1'h1:1'h1];
  assign T21656 = T18725[2'h2:2'h2];
  assign T21657 = T18725[2'h3:2'h3];
  assign T21658 = T21783 ? T21721 : T21659;
  assign T21659 = T21720 ? T21690 : T21660;
  assign T21660 = T21689 ? T21675 : T21661;
  assign T21661 = T21674 ? twiddle4_1_401_imag : twiddle4_1_400_imag;
  assign twiddle4_1_400_imag = T21664 + T21662;
  assign T21662 = $signed(T21663) / $signed(22'h100000);
  assign T21663 = $signed(31'h3c424209) * $signed(16'hffff);
  assign T21664 = {T21667, T21665};
  assign T21665 = $signed(T21666) / $signed(22'h100000);
  assign T21666 = $signed(30'h158f9a75) * $signed(16'h0);
  assign T21667 = T21665[6'h2d:6'h2d];
  assign twiddle4_1_401_imag = T21670 + T21668;
  assign T21668 = $signed(T21669) / $signed(22'h100000);
  assign T21669 = $signed(31'h3c531e88) * $signed(16'hffff);
  assign T21670 = {T21673, T21671};
  assign T21671 = $signed(T21672) / $signed(22'h100000);
  assign T21672 = $signed(30'h15604012) * $signed(16'h0);
  assign T21673 = T21671[6'h2d:6'h2d];
  assign T21674 = T18725[1'h0:1'h0];
  assign T21675 = T21688 ? twiddle4_1_403_imag : twiddle4_1_402_imag;
  assign twiddle4_1_402_imag = T21678 + T21676;
  assign T21676 = $signed(T21677) / $signed(22'h100000);
  assign T21677 = $signed(31'h3c63d5d0) * $signed(16'hffff);
  assign T21678 = {T21681, T21679};
  assign T21679 = $signed(T21680) / $signed(22'h100000);
  assign T21680 = $signed(30'h1530d880) * $signed(16'h0);
  assign T21681 = T21679[6'h2d:6'h2d];
  assign twiddle4_1_403_imag = T21684 + T21682;
  assign T21682 = $signed(T21683) / $signed(22'h100000);
  assign T21683 = $signed(31'h3c7467d8) * $signed(16'hffff);
  assign T21684 = {T21687, T21685};
  assign T21685 = $signed(T21686) / $signed(22'h100000);
  assign T21686 = $signed(30'h150163dc) * $signed(16'h0);
  assign T21687 = T21685[6'h2d:6'h2d];
  assign T21688 = T18725[1'h0:1'h0];
  assign T21689 = T18725[1'h1:1'h1];
  assign T21690 = T21719 ? T21705 : T21691;
  assign T21691 = T21704 ? twiddle4_1_405_imag : twiddle4_1_404_imag;
  assign twiddle4_1_404_imag = T21694 + T21692;
  assign T21692 = $signed(T21693) / $signed(22'h100000);
  assign T21693 = $signed(31'h3c84d496) * $signed(16'hffff);
  assign T21694 = {T21697, T21695};
  assign T21695 = $signed(T21696) / $signed(22'h100000);
  assign T21696 = $signed(30'h14d1e242) * $signed(16'h0);
  assign T21697 = T21695[6'h2d:6'h2d];
  assign twiddle4_1_405_imag = T21700 + T21698;
  assign T21698 = $signed(T21699) / $signed(22'h100000);
  assign T21699 = $signed(31'h3c951bff) * $signed(16'hffff);
  assign T21700 = {T21703, T21701};
  assign T21701 = $signed(T21702) / $signed(22'h100000);
  assign T21702 = $signed(30'h14a253d1) * $signed(16'h0);
  assign T21703 = T21701[6'h2d:6'h2d];
  assign T21704 = T18725[1'h0:1'h0];
  assign T21705 = T21718 ? twiddle4_1_407_imag : twiddle4_1_406_imag;
  assign twiddle4_1_406_imag = T21708 + T21706;
  assign T21706 = $signed(T21707) / $signed(22'h100000);
  assign T21707 = $signed(31'h3ca53e08) * $signed(16'hffff);
  assign T21708 = {T21711, T21709};
  assign T21709 = $signed(T21710) / $signed(22'h100000);
  assign T21710 = $signed(30'h1472b8a5) * $signed(16'h0);
  assign T21711 = T21709[6'h2d:6'h2d];
  assign twiddle4_1_407_imag = T21714 + T21712;
  assign T21712 = $signed(T21713) / $signed(22'h100000);
  assign T21713 = $signed(31'h3cb53aaa) * $signed(16'hffff);
  assign T21714 = {T21717, T21715};
  assign T21715 = $signed(T21716) / $signed(22'h100000);
  assign T21716 = $signed(30'h144310dc) * $signed(16'h0);
  assign T21717 = T21715[6'h2d:6'h2d];
  assign T21718 = T18725[1'h0:1'h0];
  assign T21719 = T18725[1'h1:1'h1];
  assign T21720 = T18725[2'h2:2'h2];
  assign T21721 = T21782 ? T21752 : T21722;
  assign T21722 = T21751 ? T21737 : T21723;
  assign T21723 = T21736 ? twiddle4_1_409_imag : twiddle4_1_408_imag;
  assign twiddle4_1_408_imag = T21726 + T21724;
  assign T21724 = $signed(T21725) / $signed(22'h100000);
  assign T21725 = $signed(31'h3cc511d8) * $signed(16'hffff);
  assign T21726 = {T21729, T21727};
  assign T21727 = $signed(T21728) / $signed(22'h100000);
  assign T21728 = $signed(30'h14135c94) * $signed(16'h0);
  assign T21729 = T21727[6'h2d:6'h2d];
  assign twiddle4_1_409_imag = T21732 + T21730;
  assign T21730 = $signed(T21731) / $signed(22'h100000);
  assign T21731 = $signed(31'h3cd4c38a) * $signed(16'hffff);
  assign T21732 = {T21735, T21733};
  assign T21733 = $signed(T21734) / $signed(22'h100000);
  assign T21734 = $signed(30'h13e39be9) * $signed(16'h0);
  assign T21735 = T21733[6'h2d:6'h2d];
  assign T21736 = T18725[1'h0:1'h0];
  assign T21737 = T21750 ? twiddle4_1_411_imag : twiddle4_1_410_imag;
  assign twiddle4_1_410_imag = T21740 + T21738;
  assign T21738 = $signed(T21739) / $signed(22'h100000);
  assign T21739 = $signed(31'h3ce44fb6) * $signed(16'hffff);
  assign T21740 = {T21743, T21741};
  assign T21741 = $signed(T21742) / $signed(22'h100000);
  assign T21742 = $signed(30'h13b3cefa) * $signed(16'h0);
  assign T21743 = T21741[6'h2d:6'h2d];
  assign twiddle4_1_411_imag = T21746 + T21744;
  assign T21744 = $signed(T21745) / $signed(22'h100000);
  assign T21745 = $signed(31'h3cf3b653) * $signed(16'hffff);
  assign T21746 = {T21749, T21747};
  assign T21747 = $signed(T21748) / $signed(22'h100000);
  assign T21748 = $signed(30'h1383f5e3) * $signed(16'h0);
  assign T21749 = T21747[6'h2d:6'h2d];
  assign T21750 = T18725[1'h0:1'h0];
  assign T21751 = T18725[1'h1:1'h1];
  assign T21752 = T21781 ? T21767 : T21753;
  assign T21753 = T21766 ? twiddle4_1_413_imag : twiddle4_1_412_imag;
  assign twiddle4_1_412_imag = T21756 + T21754;
  assign T21754 = $signed(T21755) / $signed(22'h100000);
  assign T21755 = $signed(31'h3d02f756) * $signed(16'hffff);
  assign T21756 = {T21759, T21757};
  assign T21757 = $signed(T21758) / $signed(22'h100000);
  assign T21758 = $signed(30'h135410c2) * $signed(16'h0);
  assign T21759 = T21757[6'h2d:6'h2d];
  assign twiddle4_1_413_imag = T21762 + T21760;
  assign T21760 = $signed(T21761) / $signed(22'h100000);
  assign T21761 = $signed(31'h3d1212b7) * $signed(16'hffff);
  assign T21762 = {T21765, T21763};
  assign T21763 = $signed(T21764) / $signed(22'h100000);
  assign T21764 = $signed(30'h13241fb6) * $signed(16'h0);
  assign T21765 = T21763[6'h2d:6'h2d];
  assign T21766 = T18725[1'h0:1'h0];
  assign T21767 = T21780 ? twiddle4_1_415_imag : twiddle4_1_414_imag;
  assign twiddle4_1_414_imag = T21770 + T21768;
  assign T21768 = $signed(T21769) / $signed(22'h100000);
  assign T21769 = $signed(31'h3d21086c) * $signed(16'hffff);
  assign T21770 = {T21773, T21771};
  assign T21771 = $signed(T21772) / $signed(22'h100000);
  assign T21772 = $signed(30'h12f422da) * $signed(16'h0);
  assign T21773 = T21771[6'h2d:6'h2d];
  assign twiddle4_1_415_imag = T21776 + T21774;
  assign T21774 = $signed(T21775) / $signed(22'h100000);
  assign T21775 = $signed(31'h3d2fd86c) * $signed(16'hffff);
  assign T21776 = {T21779, T21777};
  assign T21777 = $signed(T21778) / $signed(22'h100000);
  assign T21778 = $signed(30'h12c41a4e) * $signed(16'h0);
  assign T21779 = T21777[6'h2d:6'h2d];
  assign T21780 = T18725[1'h0:1'h0];
  assign T21781 = T18725[1'h1:1'h1];
  assign T21782 = T18725[2'h2:2'h2];
  assign T21783 = T18725[2'h3:2'h3];
  assign T21784 = T18725[3'h4:3'h4];
  assign T21785 = T22056 ? T21914 : T21786;
  assign T21786 = T21913 ? T21849 : T21787;
  assign T21787 = T21848 ? T21818 : T21788;
  assign T21788 = T21817 ? T21803 : T21789;
  assign T21789 = T21802 ? twiddle4_1_417_imag : twiddle4_1_416_imag;
  assign twiddle4_1_416_imag = T21792 + T21790;
  assign T21790 = $signed(T21791) / $signed(22'h100000);
  assign T21791 = $signed(31'h3d3e82ad) * $signed(16'hffff);
  assign T21792 = {T21795, T21793};
  assign T21793 = $signed(T21794) / $signed(22'h100000);
  assign T21794 = $signed(30'h1294062e) * $signed(16'h0);
  assign T21795 = T21793[6'h2d:6'h2d];
  assign twiddle4_1_417_imag = T21798 + T21796;
  assign T21796 = $signed(T21797) / $signed(22'h100000);
  assign T21797 = $signed(31'h3d4d0727) * $signed(16'hffff);
  assign T21798 = {T21801, T21799};
  assign T21799 = $signed(T21800) / $signed(22'h100000);
  assign T21800 = $signed(30'h1263e699) * $signed(16'h0);
  assign T21801 = T21799[6'h2d:6'h2d];
  assign T21802 = T18725[1'h0:1'h0];
  assign T21803 = T21816 ? twiddle4_1_419_imag : twiddle4_1_418_imag;
  assign twiddle4_1_418_imag = T21806 + T21804;
  assign T21804 = $signed(T21805) / $signed(22'h100000);
  assign T21805 = $signed(31'h3d5b65d1) * $signed(16'hffff);
  assign T21806 = {T21809, T21807};
  assign T21807 = $signed(T21808) / $signed(22'h100000);
  assign T21808 = $signed(30'h1233bbab) * $signed(16'h0);
  assign T21809 = T21807[6'h2d:6'h2d];
  assign twiddle4_1_419_imag = T21812 + T21810;
  assign T21810 = $signed(T21811) / $signed(22'h100000);
  assign T21811 = $signed(31'h3d699ea2) * $signed(16'hffff);
  assign T21812 = {T21815, T21813};
  assign T21813 = $signed(T21814) / $signed(22'h100000);
  assign T21814 = $signed(30'h12038583) * $signed(16'h0);
  assign T21815 = T21813[6'h2d:6'h2d];
  assign T21816 = T18725[1'h0:1'h0];
  assign T21817 = T18725[1'h1:1'h1];
  assign T21818 = T21847 ? T21833 : T21819;
  assign T21819 = T21832 ? twiddle4_1_421_imag : twiddle4_1_420_imag;
  assign twiddle4_1_420_imag = T21822 + T21820;
  assign T21820 = $signed(T21821) / $signed(22'h100000);
  assign T21821 = $signed(31'h3d77b191) * $signed(16'hffff);
  assign T21822 = {T21825, T21823};
  assign T21823 = $signed(T21824) / $signed(22'h100000);
  assign T21824 = $signed(30'h11d3443f) * $signed(16'h0);
  assign T21825 = T21823[6'h2d:6'h2d];
  assign twiddle4_1_421_imag = T21828 + T21826;
  assign T21826 = $signed(T21827) / $signed(22'h100000);
  assign T21827 = $signed(31'h3d859e96) * $signed(16'hffff);
  assign T21828 = {T21831, T21829};
  assign T21829 = $signed(T21830) / $signed(22'h100000);
  assign T21830 = $signed(30'h11a2f7fb) * $signed(16'h0);
  assign T21831 = T21829[6'h2d:6'h2d];
  assign T21832 = T18725[1'h0:1'h0];
  assign T21833 = T21846 ? twiddle4_1_423_imag : twiddle4_1_422_imag;
  assign twiddle4_1_422_imag = T21836 + T21834;
  assign T21834 = $signed(T21835) / $signed(22'h100000);
  assign T21835 = $signed(31'h3d9365a7) * $signed(16'hffff);
  assign T21836 = {T21839, T21837};
  assign T21837 = $signed(T21838) / $signed(22'h100000);
  assign T21838 = $signed(30'h1172a0d7) * $signed(16'h0);
  assign T21839 = T21837[6'h2d:6'h2d];
  assign twiddle4_1_423_imag = T21842 + T21840;
  assign T21840 = $signed(T21841) / $signed(22'h100000);
  assign T21841 = $signed(31'h3da106bd) * $signed(16'hffff);
  assign T21842 = {T21845, T21843};
  assign T21843 = $signed(T21844) / $signed(22'h100000);
  assign T21844 = $signed(30'h11423eef) * $signed(16'h0);
  assign T21845 = T21843[6'h2d:6'h2d];
  assign T21846 = T18725[1'h0:1'h0];
  assign T21847 = T18725[1'h1:1'h1];
  assign T21848 = T18725[2'h2:2'h2];
  assign T21849 = T21912 ? T21880 : T21850;
  assign T21850 = T21879 ? T21865 : T21851;
  assign T21851 = T21864 ? twiddle4_1_425_imag : twiddle4_1_424_imag;
  assign twiddle4_1_424_imag = T21854 + T21852;
  assign T21852 = $signed(T21853) / $signed(22'h100000);
  assign T21853 = $signed(31'h3dae81ce) * $signed(16'hffff);
  assign T21854 = {T21857, T21855};
  assign T21855 = $signed(T21856) / $signed(22'h100000);
  assign T21856 = $signed(30'h1111d262) * $signed(16'h0);
  assign T21857 = T21855[6'h2d:6'h2d];
  assign twiddle4_1_425_imag = T21860 + T21858;
  assign T21858 = $signed(T21859) / $signed(22'h100000);
  assign T21859 = $signed(31'h3dbbd6d4) * $signed(16'hffff);
  assign T21860 = {T21863, T21861};
  assign T21861 = $signed(T21862) / $signed(22'h100000);
  assign T21862 = $signed(30'h10e15b4e) * $signed(16'h0);
  assign T21863 = T21861[6'h2d:6'h2d];
  assign T21864 = T18725[1'h0:1'h0];
  assign T21865 = T21878 ? twiddle4_1_427_imag : twiddle4_1_426_imag;
  assign twiddle4_1_426_imag = T21868 + T21866;
  assign T21866 = $signed(T21867) / $signed(22'h100000);
  assign T21867 = $signed(31'h3dc905c4) * $signed(16'hffff);
  assign T21868 = {T21871, T21869};
  assign T21869 = $signed(T21870) / $signed(22'h100000);
  assign T21870 = $signed(30'h10b0d9cf) * $signed(16'h0);
  assign T21871 = T21869[6'h2d:6'h2d];
  assign twiddle4_1_427_imag = T21874 + T21872;
  assign T21872 = $signed(T21873) / $signed(22'h100000);
  assign T21873 = $signed(31'h3dd60e98) * $signed(16'hffff);
  assign T21874 = {T21877, T21875};
  assign T21875 = $signed(T21876) / $signed(22'h100000);
  assign T21876 = $signed(30'h10804e05) * $signed(16'h0);
  assign T21877 = T21875[6'h2d:6'h2d];
  assign T21878 = T18725[1'h0:1'h0];
  assign T21879 = T18725[1'h1:1'h1];
  assign T21880 = T21911 ? T21895 : T21881;
  assign T21881 = T21894 ? twiddle4_1_429_imag : twiddle4_1_428_imag;
  assign twiddle4_1_428_imag = T21884 + T21882;
  assign T21882 = $signed(T21883) / $signed(22'h100000);
  assign T21883 = $signed(31'h3de2f147) * $signed(16'hffff);
  assign T21884 = {T21887, T21885};
  assign T21885 = $signed(T21886) / $signed(22'h100000);
  assign T21886 = $signed(30'h104fb80e) * $signed(16'h0);
  assign T21887 = T21885[6'h2d:6'h2d];
  assign twiddle4_1_429_imag = T21890 + T21888;
  assign T21888 = $signed(T21889) / $signed(22'h100000);
  assign T21889 = $signed(31'h3defadca) * $signed(16'hffff);
  assign T21890 = {T21893, T21891};
  assign T21891 = $signed(T21892) / $signed(22'h100000);
  assign T21892 = $signed(30'h101f1806) * $signed(16'h0);
  assign T21893 = T21891[6'h2d:6'h2d];
  assign T21894 = T18725[1'h0:1'h0];
  assign T21895 = T21910 ? twiddle4_1_431_imag : twiddle4_1_430_imag;
  assign twiddle4_1_430_imag = T21898 + T21896;
  assign T21896 = $signed(T21897) / $signed(22'h100000);
  assign T21897 = $signed(31'h3dfc4418) * $signed(16'hffff);
  assign T21898 = {T21901, T21899};
  assign T21899 = $signed(T21900) / $signed(22'h100000);
  assign T21900 = $signed(29'hfee6e0d) * $signed(16'h0);
  assign T21901 = T21902 ? 2'h3 : 2'h0;
  assign T21902 = T21899[6'h2c:6'h2c];
  assign twiddle4_1_431_imag = T21905 + T21903;
  assign T21903 = $signed(T21904) / $signed(22'h100000);
  assign T21904 = $signed(31'h3e08b429) * $signed(16'hffff);
  assign T21905 = {T21908, T21906};
  assign T21906 = $signed(T21907) / $signed(22'h100000);
  assign T21907 = $signed(29'hfbdba40) * $signed(16'h0);
  assign T21908 = T21909 ? 2'h3 : 2'h0;
  assign T21909 = T21906[6'h2c:6'h2c];
  assign T21910 = T18725[1'h0:1'h0];
  assign T21911 = T18725[1'h1:1'h1];
  assign T21912 = T18725[2'h2:2'h2];
  assign T21913 = T18725[2'h3:2'h3];
  assign T21914 = T22055 ? T21985 : T21915;
  assign T21915 = T21984 ? T21950 : T21916;
  assign T21916 = T21949 ? T21933 : T21917;
  assign T21917 = T21932 ? twiddle4_1_433_imag : twiddle4_1_432_imag;
  assign twiddle4_1_432_imag = T21920 + T21918;
  assign T21918 = $signed(T21919) / $signed(22'h100000);
  assign T21919 = $signed(31'h3e14fdf7) * $signed(16'hffff);
  assign T21920 = {T21923, T21921};
  assign T21921 = $signed(T21922) / $signed(22'h100000);
  assign T21922 = $signed(29'hf8cfcbd) * $signed(16'h0);
  assign T21923 = T21924 ? 2'h3 : 2'h0;
  assign T21924 = T21921[6'h2c:6'h2c];
  assign twiddle4_1_433_imag = T21927 + T21925;
  assign T21925 = $signed(T21926) / $signed(22'h100000);
  assign T21926 = $signed(31'h3e212179) * $signed(16'hffff);
  assign T21927 = {T21930, T21928};
  assign T21928 = $signed(T21929) / $signed(22'h100000);
  assign T21929 = $signed(29'hf5c35a3) * $signed(16'h0);
  assign T21930 = T21931 ? 2'h3 : 2'h0;
  assign T21931 = T21928[6'h2c:6'h2c];
  assign T21932 = T18725[1'h0:1'h0];
  assign T21933 = T21948 ? twiddle4_1_435_imag : twiddle4_1_434_imag;
  assign twiddle4_1_434_imag = T21936 + T21934;
  assign T21934 = $signed(T21935) / $signed(22'h100000);
  assign T21935 = $signed(31'h3e2d1ea7) * $signed(16'hffff);
  assign T21936 = {T21939, T21937};
  assign T21937 = $signed(T21938) / $signed(22'h100000);
  assign T21938 = $signed(29'hf2b650f) * $signed(16'h0);
  assign T21939 = T21940 ? 2'h3 : 2'h0;
  assign T21940 = T21937[6'h2c:6'h2c];
  assign twiddle4_1_435_imag = T21943 + T21941;
  assign T21941 = $signed(T21942) / $signed(22'h100000);
  assign T21942 = $signed(31'h3e38f57c) * $signed(16'hffff);
  assign T21943 = {T21946, T21944};
  assign T21944 = $signed(T21945) / $signed(22'h100000);
  assign T21945 = $signed(29'hefa8b1f) * $signed(16'h0);
  assign T21946 = T21947 ? 2'h3 : 2'h0;
  assign T21947 = T21944[6'h2c:6'h2c];
  assign T21948 = T18725[1'h0:1'h0];
  assign T21949 = T18725[1'h1:1'h1];
  assign T21950 = T21983 ? T21967 : T21951;
  assign T21951 = T21966 ? twiddle4_1_437_imag : twiddle4_1_436_imag;
  assign twiddle4_1_436_imag = T21954 + T21952;
  assign T21952 = $signed(T21953) / $signed(22'h100000);
  assign T21953 = $signed(31'h3e44a5ee) * $signed(16'hffff);
  assign T21954 = {T21957, T21955};
  assign T21955 = $signed(T21956) / $signed(22'h100000);
  assign T21956 = $signed(29'hec9a7f2) * $signed(16'h0);
  assign T21957 = T21958 ? 2'h3 : 2'h0;
  assign T21958 = T21955[6'h2c:6'h2c];
  assign twiddle4_1_437_imag = T21961 + T21959;
  assign T21959 = $signed(T21960) / $signed(22'h100000);
  assign T21960 = $signed(31'h3e502ff8) * $signed(16'hffff);
  assign T21961 = {T21964, T21962};
  assign T21962 = $signed(T21963) / $signed(22'h100000);
  assign T21963 = $signed(29'he98bba6) * $signed(16'h0);
  assign T21964 = T21965 ? 2'h3 : 2'h0;
  assign T21965 = T21962[6'h2c:6'h2c];
  assign T21966 = T18725[1'h0:1'h0];
  assign T21967 = T21982 ? twiddle4_1_439_imag : twiddle4_1_438_imag;
  assign twiddle4_1_438_imag = T21970 + T21968;
  assign T21968 = $signed(T21969) / $signed(22'h100000);
  assign T21969 = $signed(31'h3e5b9392) * $signed(16'hffff);
  assign T21970 = {T21973, T21971};
  assign T21971 = $signed(T21972) / $signed(22'h100000);
  assign T21972 = $signed(29'he67c659) * $signed(16'h0);
  assign T21973 = T21974 ? 2'h3 : 2'h0;
  assign T21974 = T21971[6'h2c:6'h2c];
  assign twiddle4_1_439_imag = T21977 + T21975;
  assign T21975 = $signed(T21976) / $signed(22'h100000);
  assign T21976 = $signed(31'h3e66d0b4) * $signed(16'hffff);
  assign T21977 = {T21980, T21978};
  assign T21978 = $signed(T21979) / $signed(22'h100000);
  assign T21979 = $signed(29'he36c829) * $signed(16'h0);
  assign T21980 = T21981 ? 2'h3 : 2'h0;
  assign T21981 = T21978[6'h2c:6'h2c];
  assign T21982 = T18725[1'h0:1'h0];
  assign T21983 = T18725[1'h1:1'h1];
  assign T21984 = T18725[2'h2:2'h2];
  assign T21985 = T22054 ? T22020 : T21986;
  assign T21986 = T22019 ? T22003 : T21987;
  assign T21987 = T22002 ? twiddle4_1_441_imag : twiddle4_1_440_imag;
  assign twiddle4_1_440_imag = T21990 + T21988;
  assign T21988 = $signed(T21989) / $signed(22'h100000);
  assign T21989 = $signed(31'h3e71e758) * $signed(16'hffff);
  assign T21990 = {T21993, T21991};
  assign T21991 = $signed(T21992) / $signed(22'h100000);
  assign T21992 = $signed(29'he05c135) * $signed(16'h0);
  assign T21993 = T21994 ? 2'h3 : 2'h0;
  assign T21994 = T21991[6'h2c:6'h2c];
  assign twiddle4_1_441_imag = T21997 + T21995;
  assign T21995 = $signed(T21996) / $signed(22'h100000);
  assign T21996 = $signed(31'h3e7cd778) * $signed(16'hffff);
  assign T21997 = {T22000, T21998};
  assign T21998 = $signed(T21999) / $signed(22'h100000);
  assign T21999 = $signed(29'hdd4b19a) * $signed(16'h0);
  assign T22000 = T22001 ? 2'h3 : 2'h0;
  assign T22001 = T21998[6'h2c:6'h2c];
  assign T22002 = T18725[1'h0:1'h0];
  assign T22003 = T22018 ? twiddle4_1_443_imag : twiddle4_1_442_imag;
  assign twiddle4_1_442_imag = T22006 + T22004;
  assign T22004 = $signed(T22005) / $signed(22'h100000);
  assign T22005 = $signed(31'h3e87a10b) * $signed(16'hffff);
  assign T22006 = {T22009, T22007};
  assign T22007 = $signed(T22008) / $signed(22'h100000);
  assign T22008 = $signed(29'hda39977) * $signed(16'h0);
  assign T22009 = T22010 ? 2'h3 : 2'h0;
  assign T22010 = T22007[6'h2c:6'h2c];
  assign twiddle4_1_443_imag = T22013 + T22011;
  assign T22011 = $signed(T22012) / $signed(22'h100000);
  assign T22012 = $signed(31'h3e92440d) * $signed(16'hffff);
  assign T22013 = {T22016, T22014};
  assign T22014 = $signed(T22015) / $signed(22'h100000);
  assign T22015 = $signed(29'hd7278ea) * $signed(16'h0);
  assign T22016 = T22017 ? 2'h3 : 2'h0;
  assign T22017 = T22014[6'h2c:6'h2c];
  assign T22018 = T18725[1'h0:1'h0];
  assign T22019 = T18725[1'h1:1'h1];
  assign T22020 = T22053 ? T22037 : T22021;
  assign T22021 = T22036 ? twiddle4_1_445_imag : twiddle4_1_444_imag;
  assign twiddle4_1_444_imag = T22024 + T22022;
  assign T22022 = $signed(T22023) / $signed(22'h100000);
  assign T22023 = $signed(31'h3e9cc076) * $signed(16'hffff);
  assign T22024 = {T22027, T22025};
  assign T22025 = $signed(T22026) / $signed(22'h100000);
  assign T22026 = $signed(29'hd415012) * $signed(16'h0);
  assign T22027 = T22028 ? 2'h3 : 2'h0;
  assign T22028 = T22025[6'h2c:6'h2c];
  assign twiddle4_1_445_imag = T22031 + T22029;
  assign T22029 = $signed(T22030) / $signed(22'h100000);
  assign T22030 = $signed(31'h3ea7163f) * $signed(16'hffff);
  assign T22031 = {T22034, T22032};
  assign T22032 = $signed(T22033) / $signed(22'h100000);
  assign T22033 = $signed(29'hd101f0d) * $signed(16'h0);
  assign T22034 = T22035 ? 2'h3 : 2'h0;
  assign T22035 = T22032[6'h2c:6'h2c];
  assign T22036 = T18725[1'h0:1'h0];
  assign T22037 = T22052 ? twiddle4_1_447_imag : twiddle4_1_446_imag;
  assign twiddle4_1_446_imag = T22040 + T22038;
  assign T22038 = $signed(T22039) / $signed(22'h100000);
  assign T22039 = $signed(31'h3eb14562) * $signed(16'hffff);
  assign T22040 = {T22043, T22041};
  assign T22041 = $signed(T22042) / $signed(22'h100000);
  assign T22042 = $signed(29'hcdee5f9) * $signed(16'h0);
  assign T22043 = T22044 ? 2'h3 : 2'h0;
  assign T22044 = T22041[6'h2c:6'h2c];
  assign twiddle4_1_447_imag = T22047 + T22045;
  assign T22045 = $signed(T22046) / $signed(22'h100000);
  assign T22046 = $signed(31'h3ebb4dda) * $signed(16'hffff);
  assign T22047 = {T22050, T22048};
  assign T22048 = $signed(T22049) / $signed(22'h100000);
  assign T22049 = $signed(29'hcada4f4) * $signed(16'h0);
  assign T22050 = T22051 ? 2'h3 : 2'h0;
  assign T22051 = T22048[6'h2c:6'h2c];
  assign T22052 = T18725[1'h0:1'h0];
  assign T22053 = T18725[1'h1:1'h1];
  assign T22054 = T18725[2'h2:2'h2];
  assign T22055 = T18725[2'h3:2'h3];
  assign T22056 = T18725[3'h4:3'h4];
  assign T22057 = T18725[3'h5:3'h5];
  assign T22058 = T22631 ? T22345 : T22059;
  assign T22059 = T22344 ? T22202 : T22060;
  assign T22060 = T22201 ? T22131 : T22061;
  assign T22061 = T22130 ? T22096 : T22062;
  assign T22062 = T22095 ? T22079 : T22063;
  assign T22063 = T22078 ? twiddle4_1_449_imag : twiddle4_1_448_imag;
  assign twiddle4_1_448_imag = T22066 + T22064;
  assign T22064 = $signed(T22065) / $signed(22'h100000);
  assign T22065 = $signed(31'h3ec52f9f) * $signed(16'hffff);
  assign T22066 = {T22069, T22067};
  assign T22067 = $signed(T22068) / $signed(22'h100000);
  assign T22068 = $signed(29'hc7c5c1e) * $signed(16'h0);
  assign T22069 = T22070 ? 2'h3 : 2'h0;
  assign T22070 = T22067[6'h2c:6'h2c];
  assign twiddle4_1_449_imag = T22073 + T22071;
  assign T22071 = $signed(T22072) / $signed(22'h100000);
  assign T22072 = $signed(31'h3eceeaad) * $signed(16'hffff);
  assign T22073 = {T22076, T22074};
  assign T22074 = $signed(T22075) / $signed(22'h100000);
  assign T22075 = $signed(29'hc4b0b93) * $signed(16'h0);
  assign T22076 = T22077 ? 2'h3 : 2'h0;
  assign T22077 = T22074[6'h2c:6'h2c];
  assign T22078 = T18725[1'h0:1'h0];
  assign T22079 = T22094 ? twiddle4_1_451_imag : twiddle4_1_450_imag;
  assign twiddle4_1_450_imag = T22082 + T22080;
  assign T22080 = $signed(T22081) / $signed(22'h100000);
  assign T22081 = $signed(31'h3ed87efb) * $signed(16'hffff);
  assign T22082 = {T22085, T22083};
  assign T22083 = $signed(T22084) / $signed(22'h100000);
  assign T22084 = $signed(29'hc19b374) * $signed(16'h0);
  assign T22085 = T22086 ? 2'h3 : 2'h0;
  assign T22086 = T22083[6'h2c:6'h2c];
  assign twiddle4_1_451_imag = T22089 + T22087;
  assign T22087 = $signed(T22088) / $signed(22'h100000);
  assign T22088 = $signed(31'h3ee1ec86) * $signed(16'hffff);
  assign T22089 = {T22092, T22090};
  assign T22090 = $signed(T22091) / $signed(22'h100000);
  assign T22091 = $signed(29'hbe853dd) * $signed(16'h0);
  assign T22092 = T22093 ? 2'h3 : 2'h0;
  assign T22093 = T22090[6'h2c:6'h2c];
  assign T22094 = T18725[1'h0:1'h0];
  assign T22095 = T18725[1'h1:1'h1];
  assign T22096 = T22129 ? T22113 : T22097;
  assign T22097 = T22112 ? twiddle4_1_453_imag : twiddle4_1_452_imag;
  assign twiddle4_1_452_imag = T22100 + T22098;
  assign T22098 = $signed(T22099) / $signed(22'h100000);
  assign T22099 = $signed(31'h3eeb3347) * $signed(16'hffff);
  assign T22100 = {T22103, T22101};
  assign T22101 = $signed(T22102) / $signed(22'h100000);
  assign T22102 = $signed(29'hbb6ecef) * $signed(16'h0);
  assign T22103 = T22104 ? 2'h3 : 2'h0;
  assign T22104 = T22101[6'h2c:6'h2c];
  assign twiddle4_1_453_imag = T22107 + T22105;
  assign T22105 = $signed(T22106) / $signed(22'h100000);
  assign T22106 = $signed(31'h3ef45338) * $signed(16'hffff);
  assign T22107 = {T22110, T22108};
  assign T22108 = $signed(T22109) / $signed(22'h100000);
  assign T22109 = $signed(29'hb857ec6) * $signed(16'h0);
  assign T22110 = T22111 ? 2'h3 : 2'h0;
  assign T22111 = T22108[6'h2c:6'h2c];
  assign T22112 = T18725[1'h0:1'h0];
  assign T22113 = T22128 ? twiddle4_1_455_imag : twiddle4_1_454_imag;
  assign twiddle4_1_454_imag = T22116 + T22114;
  assign T22114 = $signed(T22115) / $signed(22'h100000);
  assign T22115 = $signed(31'h3efd4c53) * $signed(16'hffff);
  assign T22116 = {T22119, T22117};
  assign T22117 = $signed(T22118) / $signed(22'h100000);
  assign T22118 = $signed(29'hb540982) * $signed(16'h0);
  assign T22119 = T22120 ? 2'h3 : 2'h0;
  assign T22120 = T22117[6'h2c:6'h2c];
  assign twiddle4_1_455_imag = T22123 + T22121;
  assign T22121 = $signed(T22122) / $signed(22'h100000);
  assign T22122 = $signed(31'h3f061e94) * $signed(16'hffff);
  assign T22123 = {T22126, T22124};
  assign T22124 = $signed(T22125) / $signed(22'h100000);
  assign T22125 = $signed(29'hb228d41) * $signed(16'h0);
  assign T22126 = T22127 ? 2'h3 : 2'h0;
  assign T22127 = T22124[6'h2c:6'h2c];
  assign T22128 = T18725[1'h0:1'h0];
  assign T22129 = T18725[1'h1:1'h1];
  assign T22130 = T18725[2'h2:2'h2];
  assign T22131 = T22200 ? T22166 : T22132;
  assign T22132 = T22165 ? T22149 : T22133;
  assign T22133 = T22148 ? twiddle4_1_457_imag : twiddle4_1_456_imag;
  assign twiddle4_1_456_imag = T22136 + T22134;
  assign T22134 = $signed(T22135) / $signed(22'h100000);
  assign T22135 = $signed(31'h3f0ec9f4) * $signed(16'hffff);
  assign T22136 = {T22139, T22137};
  assign T22137 = $signed(T22138) / $signed(22'h100000);
  assign T22138 = $signed(29'haf10a22) * $signed(16'h0);
  assign T22139 = T22140 ? 2'h3 : 2'h0;
  assign T22140 = T22137[6'h2c:6'h2c];
  assign twiddle4_1_457_imag = T22143 + T22141;
  assign T22141 = $signed(T22142) / $signed(22'h100000);
  assign T22142 = $signed(31'h3f174e6f) * $signed(16'hffff);
  assign T22143 = {T22146, T22144};
  assign T22144 = $signed(T22145) / $signed(22'h100000);
  assign T22145 = $signed(29'habf8043) * $signed(16'h0);
  assign T22146 = T22147 ? 2'h3 : 2'h0;
  assign T22147 = T22144[6'h2c:6'h2c];
  assign T22148 = T18725[1'h0:1'h0];
  assign T22149 = T22164 ? twiddle4_1_459_imag : twiddle4_1_458_imag;
  assign twiddle4_1_458_imag = T22152 + T22150;
  assign T22150 = $signed(T22151) / $signed(22'h100000);
  assign T22151 = $signed(31'h3f1fabff) * $signed(16'hffff);
  assign T22152 = {T22155, T22153};
  assign T22153 = $signed(T22154) / $signed(22'h100000);
  assign T22154 = $signed(29'ha8defc2) * $signed(16'h0);
  assign T22155 = T22156 ? 2'h3 : 2'h0;
  assign T22156 = T22153[6'h2c:6'h2c];
  assign twiddle4_1_459_imag = T22159 + T22157;
  assign T22157 = $signed(T22158) / $signed(22'h100000);
  assign T22158 = $signed(31'h3f27e29f) * $signed(16'hffff);
  assign T22159 = {T22162, T22160};
  assign T22160 = $signed(T22161) / $signed(22'h100000);
  assign T22161 = $signed(29'ha5c58bf) * $signed(16'h0);
  assign T22162 = T22163 ? 2'h3 : 2'h0;
  assign T22163 = T22160[6'h2c:6'h2c];
  assign T22164 = T18725[1'h0:1'h0];
  assign T22165 = T18725[1'h1:1'h1];
  assign T22166 = T22199 ? T22183 : T22167;
  assign T22167 = T22182 ? twiddle4_1_461_imag : twiddle4_1_460_imag;
  assign twiddle4_1_460_imag = T22170 + T22168;
  assign T22168 = $signed(T22169) / $signed(22'h100000);
  assign T22169 = $signed(31'h3f2ff249) * $signed(16'hffff);
  assign T22170 = {T22173, T22171};
  assign T22171 = $signed(T22172) / $signed(22'h100000);
  assign T22172 = $signed(29'ha2abb58) * $signed(16'h0);
  assign T22173 = T22174 ? 2'h3 : 2'h0;
  assign T22174 = T22171[6'h2c:6'h2c];
  assign twiddle4_1_461_imag = T22177 + T22175;
  assign T22175 = $signed(T22176) / $signed(22'h100000);
  assign T22176 = $signed(31'h3f37daf9) * $signed(16'hffff);
  assign T22177 = {T22180, T22178};
  assign T22178 = $signed(T22179) / $signed(22'h100000);
  assign T22179 = $signed(29'h9f917ab) * $signed(16'h0);
  assign T22180 = T22181 ? 2'h3 : 2'h0;
  assign T22181 = T22178[6'h2c:6'h2c];
  assign T22182 = T18725[1'h0:1'h0];
  assign T22183 = T22198 ? twiddle4_1_463_imag : twiddle4_1_462_imag;
  assign twiddle4_1_462_imag = T22186 + T22184;
  assign T22184 = $signed(T22185) / $signed(22'h100000);
  assign T22185 = $signed(31'h3f3f9cab) * $signed(16'hffff);
  assign T22186 = {T22189, T22187};
  assign T22187 = $signed(T22188) / $signed(22'h100000);
  assign T22188 = $signed(29'h9c76dd8) * $signed(16'h0);
  assign T22189 = T22190 ? 2'h3 : 2'h0;
  assign T22190 = T22187[6'h2c:6'h2c];
  assign twiddle4_1_463_imag = T22193 + T22191;
  assign T22191 = $signed(T22192) / $signed(22'h100000);
  assign T22192 = $signed(31'h3f473758) * $signed(16'hffff);
  assign T22193 = {T22196, T22194};
  assign T22194 = $signed(T22195) / $signed(22'h100000);
  assign T22195 = $signed(29'h995bdfc) * $signed(16'h0);
  assign T22196 = T22197 ? 2'h3 : 2'h0;
  assign T22197 = T22194[6'h2c:6'h2c];
  assign T22198 = T18725[1'h0:1'h0];
  assign T22199 = T18725[1'h1:1'h1];
  assign T22200 = T18725[2'h2:2'h2];
  assign T22201 = T18725[2'h3:2'h3];
  assign T22202 = T22343 ? T22273 : T22203;
  assign T22203 = T22272 ? T22238 : T22204;
  assign T22204 = T22237 ? T22221 : T22205;
  assign T22205 = T22220 ? twiddle4_1_465_imag : twiddle4_1_464_imag;
  assign twiddle4_1_464_imag = T22208 + T22206;
  assign T22206 = $signed(T22207) / $signed(22'h100000);
  assign T22207 = $signed(31'h3f4eaafe) * $signed(16'hffff);
  assign T22208 = {T22211, T22209};
  assign T22209 = $signed(T22210) / $signed(22'h100000);
  assign T22210 = $signed(29'h9640837) * $signed(16'h0);
  assign T22211 = T22212 ? 2'h3 : 2'h0;
  assign T22212 = T22209[6'h2c:6'h2c];
  assign twiddle4_1_465_imag = T22215 + T22213;
  assign T22213 = $signed(T22214) / $signed(22'h100000);
  assign T22214 = $signed(31'h3f55f796) * $signed(16'hffff);
  assign T22215 = {T22218, T22216};
  assign T22216 = $signed(T22217) / $signed(22'h100000);
  assign T22217 = $signed(29'h9324ca6) * $signed(16'h0);
  assign T22218 = T22219 ? 2'h3 : 2'h0;
  assign T22219 = T22216[6'h2c:6'h2c];
  assign T22220 = T18725[1'h0:1'h0];
  assign T22221 = T22236 ? twiddle4_1_467_imag : twiddle4_1_466_imag;
  assign twiddle4_1_466_imag = T22224 + T22222;
  assign T22222 = $signed(T22223) / $signed(22'h100000);
  assign T22223 = $signed(31'h3f5d1d1c) * $signed(16'hffff);
  assign T22224 = {T22227, T22225};
  assign T22225 = $signed(T22226) / $signed(22'h100000);
  assign T22226 = $signed(29'h9008b6a) * $signed(16'h0);
  assign T22227 = T22228 ? 2'h3 : 2'h0;
  assign T22228 = T22225[6'h2c:6'h2c];
  assign twiddle4_1_467_imag = T22231 + T22229;
  assign T22229 = $signed(T22230) / $signed(22'h100000);
  assign T22230 = $signed(31'h3f641b8d) * $signed(16'hffff);
  assign T22231 = {T22234, T22232};
  assign T22232 = $signed(T22233) / $signed(22'h100000);
  assign T22233 = $signed(29'h8cec4a0) * $signed(16'h0);
  assign T22234 = T22235 ? 2'h3 : 2'h0;
  assign T22235 = T22232[6'h2c:6'h2c];
  assign T22236 = T18725[1'h0:1'h0];
  assign T22237 = T18725[1'h1:1'h1];
  assign T22238 = T22271 ? T22255 : T22239;
  assign T22239 = T22254 ? twiddle4_1_469_imag : twiddle4_1_468_imag;
  assign twiddle4_1_468_imag = T22242 + T22240;
  assign T22240 = $signed(T22241) / $signed(22'h100000);
  assign T22241 = $signed(31'h3f6af2e3) * $signed(16'hffff);
  assign T22242 = {T22245, T22243};
  assign T22243 = $signed(T22244) / $signed(22'h100000);
  assign T22244 = $signed(29'h89cf867) * $signed(16'h0);
  assign T22245 = T22246 ? 2'h3 : 2'h0;
  assign T22246 = T22243[6'h2c:6'h2c];
  assign twiddle4_1_469_imag = T22249 + T22247;
  assign T22247 = $signed(T22248) / $signed(22'h100000);
  assign T22248 = $signed(31'h3f71a31a) * $signed(16'hffff);
  assign T22249 = {T22252, T22250};
  assign T22250 = $signed(T22251) / $signed(22'h100000);
  assign T22251 = $signed(29'h86b26de) * $signed(16'h0);
  assign T22252 = T22253 ? 2'h3 : 2'h0;
  assign T22253 = T22250[6'h2c:6'h2c];
  assign T22254 = T18725[1'h0:1'h0];
  assign T22255 = T22270 ? twiddle4_1_471_imag : twiddle4_1_470_imag;
  assign twiddle4_1_470_imag = T22258 + T22256;
  assign T22256 = $signed(T22257) / $signed(22'h100000);
  assign T22257 = $signed(31'h3f782c2f) * $signed(16'hffff);
  assign T22258 = {T22261, T22259};
  assign T22259 = $signed(T22260) / $signed(22'h100000);
  assign T22260 = $signed(29'h8395023) * $signed(16'h0);
  assign T22261 = T22262 ? 2'h3 : 2'h0;
  assign T22262 = T22259[6'h2c:6'h2c];
  assign twiddle4_1_471_imag = T22265 + T22263;
  assign T22263 = $signed(T22264) / $signed(22'h100000);
  assign T22264 = $signed(31'h3f7e8e1e) * $signed(16'hffff);
  assign T22265 = {T22268, T22266};
  assign T22266 = $signed(T22267) / $signed(22'h100000);
  assign T22267 = $signed(29'h8077456) * $signed(16'h0);
  assign T22268 = T22269 ? 2'h3 : 2'h0;
  assign T22269 = T22266[6'h2c:6'h2c];
  assign T22270 = T18725[1'h0:1'h0];
  assign T22271 = T18725[1'h1:1'h1];
  assign T22272 = T18725[2'h2:2'h2];
  assign T22273 = T22342 ? T22308 : T22274;
  assign T22274 = T22307 ? T22291 : T22275;
  assign T22275 = T22290 ? twiddle4_1_473_imag : twiddle4_1_472_imag;
  assign twiddle4_1_472_imag = T22278 + T22276;
  assign T22276 = $signed(T22277) / $signed(22'h100000);
  assign T22277 = $signed(31'h3f84c8e1) * $signed(16'hffff);
  assign T22278 = {T22281, T22279};
  assign T22279 = $signed(T22280) / $signed(22'h100000);
  assign T22280 = $signed(28'h7d59395) * $signed(16'h0);
  assign T22281 = T22282 ? 3'h7 : 3'h0;
  assign T22282 = T22279[6'h2b:6'h2b];
  assign twiddle4_1_473_imag = T22285 + T22283;
  assign T22283 = $signed(T22284) / $signed(22'h100000);
  assign T22284 = $signed(31'h3f8adc76) * $signed(16'hffff);
  assign T22285 = {T22288, T22286};
  assign T22286 = $signed(T22287) / $signed(22'h100000);
  assign T22287 = $signed(28'h7a3adff) * $signed(16'h0);
  assign T22288 = T22289 ? 3'h7 : 3'h0;
  assign T22289 = T22286[6'h2b:6'h2b];
  assign T22290 = T18725[1'h0:1'h0];
  assign T22291 = T22306 ? twiddle4_1_475_imag : twiddle4_1_474_imag;
  assign twiddle4_1_474_imag = T22294 + T22292;
  assign T22292 = $signed(T22293) / $signed(22'h100000);
  assign T22293 = $signed(31'h3f90c8d9) * $signed(16'hffff);
  assign T22294 = {T22297, T22295};
  assign T22295 = $signed(T22296) / $signed(22'h100000);
  assign T22296 = $signed(28'h771c3b2) * $signed(16'h0);
  assign T22297 = T22298 ? 3'h7 : 3'h0;
  assign T22298 = T22295[6'h2b:6'h2b];
  assign twiddle4_1_475_imag = T22301 + T22299;
  assign T22299 = $signed(T22300) / $signed(22'h100000);
  assign T22300 = $signed(31'h3f968e07) * $signed(16'hffff);
  assign T22301 = {T22304, T22302};
  assign T22302 = $signed(T22303) / $signed(22'h100000);
  assign T22303 = $signed(28'h73fd4ce) * $signed(16'h0);
  assign T22304 = T22305 ? 3'h7 : 3'h0;
  assign T22305 = T22302[6'h2b:6'h2b];
  assign T22306 = T18725[1'h0:1'h0];
  assign T22307 = T18725[1'h1:1'h1];
  assign T22308 = T22341 ? T22325 : T22309;
  assign T22309 = T22324 ? twiddle4_1_477_imag : twiddle4_1_476_imag;
  assign twiddle4_1_476_imag = T22312 + T22310;
  assign T22310 = $signed(T22311) / $signed(22'h100000);
  assign T22311 = $signed(31'h3f9c2bfa) * $signed(16'hffff);
  assign T22312 = {T22315, T22313};
  assign T22313 = $signed(T22314) / $signed(22'h100000);
  assign T22314 = $signed(28'h70de171) * $signed(16'h0);
  assign T22315 = T22316 ? 3'h7 : 3'h0;
  assign T22316 = T22313[6'h2b:6'h2b];
  assign twiddle4_1_477_imag = T22319 + T22317;
  assign T22317 = $signed(T22318) / $signed(22'h100000);
  assign T22318 = $signed(31'h3fa1a2b1) * $signed(16'hffff);
  assign T22319 = {T22322, T22320};
  assign T22320 = $signed(T22321) / $signed(22'h100000);
  assign T22321 = $signed(28'h6dbe9bb) * $signed(16'h0);
  assign T22322 = T22323 ? 3'h7 : 3'h0;
  assign T22323 = T22320[6'h2b:6'h2b];
  assign T22324 = T18725[1'h0:1'h0];
  assign T22325 = T22340 ? twiddle4_1_479_imag : twiddle4_1_478_imag;
  assign twiddle4_1_478_imag = T22328 + T22326;
  assign T22326 = $signed(T22327) / $signed(22'h100000);
  assign T22327 = $signed(31'h3fa6f228) * $signed(16'hffff);
  assign T22328 = {T22331, T22329};
  assign T22329 = $signed(T22330) / $signed(22'h100000);
  assign T22330 = $signed(28'h6a9edc9) * $signed(16'h0);
  assign T22331 = T22332 ? 3'h7 : 3'h0;
  assign T22332 = T22329[6'h2b:6'h2b];
  assign twiddle4_1_479_imag = T22335 + T22333;
  assign T22333 = $signed(T22334) / $signed(22'h100000);
  assign T22334 = $signed(31'h3fac1a5b) * $signed(16'hffff);
  assign T22335 = {T22338, T22336};
  assign T22336 = $signed(T22337) / $signed(22'h100000);
  assign T22337 = $signed(28'h677edba) * $signed(16'h0);
  assign T22338 = T22339 ? 3'h7 : 3'h0;
  assign T22339 = T22336[6'h2b:6'h2b];
  assign T22340 = T18725[1'h0:1'h0];
  assign T22341 = T18725[1'h1:1'h1];
  assign T22342 = T18725[2'h2:2'h2];
  assign T22343 = T18725[2'h3:2'h3];
  assign T22344 = T18725[3'h4:3'h4];
  assign T22345 = T22630 ? T22488 : T22346;
  assign T22346 = T22487 ? T22417 : T22347;
  assign T22347 = T22416 ? T22382 : T22348;
  assign T22348 = T22381 ? T22365 : T22349;
  assign T22349 = T22364 ? twiddle4_1_481_imag : twiddle4_1_480_imag;
  assign twiddle4_1_480_imag = T22352 + T22350;
  assign T22350 = $signed(T22351) / $signed(22'h100000);
  assign T22351 = $signed(31'h3fb11b47) * $signed(16'hffff);
  assign T22352 = {T22355, T22353};
  assign T22353 = $signed(T22354) / $signed(22'h100000);
  assign T22354 = $signed(28'h645e9af) * $signed(16'h0);
  assign T22355 = T22356 ? 3'h7 : 3'h0;
  assign T22356 = T22353[6'h2b:6'h2b];
  assign twiddle4_1_481_imag = T22359 + T22357;
  assign T22357 = $signed(T22358) / $signed(22'h100000);
  assign T22358 = $signed(31'h3fb5f4ea) * $signed(16'hffff);
  assign T22359 = {T22362, T22360};
  assign T22360 = $signed(T22361) / $signed(22'h100000);
  assign T22361 = $signed(28'h613e1c4) * $signed(16'h0);
  assign T22362 = T22363 ? 3'h7 : 3'h0;
  assign T22363 = T22360[6'h2b:6'h2b];
  assign T22364 = T18725[1'h0:1'h0];
  assign T22365 = T22380 ? twiddle4_1_483_imag : twiddle4_1_482_imag;
  assign twiddle4_1_482_imag = T22368 + T22366;
  assign T22366 = $signed(T22367) / $signed(22'h100000);
  assign T22367 = $signed(31'h3fbaa73f) * $signed(16'hffff);
  assign T22368 = {T22371, T22369};
  assign T22369 = $signed(T22370) / $signed(22'h100000);
  assign T22370 = $signed(28'h5e1d61a) * $signed(16'h0);
  assign T22371 = T22372 ? 3'h7 : 3'h0;
  assign T22372 = T22369[6'h2b:6'h2b];
  assign twiddle4_1_483_imag = T22375 + T22373;
  assign T22373 = $signed(T22374) / $signed(22'h100000);
  assign T22374 = $signed(31'h3fbf3245) * $signed(16'hffff);
  assign T22375 = {T22378, T22376};
  assign T22376 = $signed(T22377) / $signed(22'h100000);
  assign T22377 = $signed(28'h5afc6cf) * $signed(16'h0);
  assign T22378 = T22379 ? 3'h7 : 3'h0;
  assign T22379 = T22376[6'h2b:6'h2b];
  assign T22380 = T18725[1'h0:1'h0];
  assign T22381 = T18725[1'h1:1'h1];
  assign T22382 = T22415 ? T22399 : T22383;
  assign T22383 = T22398 ? twiddle4_1_485_imag : twiddle4_1_484_imag;
  assign twiddle4_1_484_imag = T22386 + T22384;
  assign T22384 = $signed(T22385) / $signed(22'h100000);
  assign T22385 = $signed(31'h3fc395f9) * $signed(16'hffff);
  assign T22386 = {T22389, T22387};
  assign T22387 = $signed(T22388) / $signed(22'h100000);
  assign T22388 = $signed(28'h57db402) * $signed(16'h0);
  assign T22389 = T22390 ? 3'h7 : 3'h0;
  assign T22390 = T22387[6'h2b:6'h2b];
  assign twiddle4_1_485_imag = T22393 + T22391;
  assign T22391 = $signed(T22392) / $signed(22'h100000);
  assign T22392 = $signed(31'h3fc7d257) * $signed(16'hffff);
  assign T22393 = {T22396, T22394};
  assign T22394 = $signed(T22395) / $signed(22'h100000);
  assign T22395 = $signed(28'h54b9dd2) * $signed(16'h0);
  assign T22396 = T22397 ? 3'h7 : 3'h0;
  assign T22397 = T22394[6'h2b:6'h2b];
  assign T22398 = T18725[1'h0:1'h0];
  assign T22399 = T22414 ? twiddle4_1_487_imag : twiddle4_1_486_imag;
  assign twiddle4_1_486_imag = T22402 + T22400;
  assign T22400 = $signed(T22401) / $signed(22'h100000);
  assign T22401 = $signed(31'h3fcbe75e) * $signed(16'hffff);
  assign T22402 = {T22405, T22403};
  assign T22403 = $signed(T22404) / $signed(22'h100000);
  assign T22404 = $signed(28'h519845e) * $signed(16'h0);
  assign T22405 = T22406 ? 3'h7 : 3'h0;
  assign T22406 = T22403[6'h2b:6'h2b];
  assign twiddle4_1_487_imag = T22409 + T22407;
  assign T22407 = $signed(T22408) / $signed(22'h100000);
  assign T22408 = $signed(31'h3fcfd50a) * $signed(16'hffff);
  assign T22409 = {T22412, T22410};
  assign T22410 = $signed(T22411) / $signed(22'h100000);
  assign T22411 = $signed(28'h4e767c4) * $signed(16'h0);
  assign T22412 = T22413 ? 3'h7 : 3'h0;
  assign T22413 = T22410[6'h2b:6'h2b];
  assign T22414 = T18725[1'h0:1'h0];
  assign T22415 = T18725[1'h1:1'h1];
  assign T22416 = T18725[2'h2:2'h2];
  assign T22417 = T22486 ? T22452 : T22418;
  assign T22418 = T22451 ? T22435 : T22419;
  assign T22419 = T22434 ? twiddle4_1_489_imag : twiddle4_1_488_imag;
  assign twiddle4_1_488_imag = T22422 + T22420;
  assign T22420 = $signed(T22421) / $signed(22'h100000);
  assign T22421 = $signed(31'h3fd39b5a) * $signed(16'hffff);
  assign T22422 = {T22425, T22423};
  assign T22423 = $signed(T22424) / $signed(22'h100000);
  assign T22424 = $signed(28'h4b54824) * $signed(16'h0);
  assign T22425 = T22426 ? 3'h7 : 3'h0;
  assign T22426 = T22423[6'h2b:6'h2b];
  assign twiddle4_1_489_imag = T22429 + T22427;
  assign T22427 = $signed(T22428) / $signed(22'h100000);
  assign T22428 = $signed(31'h3fd73a4a) * $signed(16'hffff);
  assign T22429 = {T22432, T22430};
  assign T22430 = $signed(T22431) / $signed(22'h100000);
  assign T22431 = $signed(28'h483259d) * $signed(16'h0);
  assign T22432 = T22433 ? 3'h7 : 3'h0;
  assign T22433 = T22430[6'h2b:6'h2b];
  assign T22434 = T18725[1'h0:1'h0];
  assign T22435 = T22450 ? twiddle4_1_491_imag : twiddle4_1_490_imag;
  assign twiddle4_1_490_imag = T22438 + T22436;
  assign T22436 = $signed(T22437) / $signed(22'h100000);
  assign T22437 = $signed(31'h3fdab1d9) * $signed(16'hffff);
  assign T22438 = {T22441, T22439};
  assign T22439 = $signed(T22440) / $signed(22'h100000);
  assign T22440 = $signed(28'h451004d) * $signed(16'h0);
  assign T22441 = T22442 ? 3'h7 : 3'h0;
  assign T22442 = T22439[6'h2b:6'h2b];
  assign twiddle4_1_491_imag = T22445 + T22443;
  assign T22443 = $signed(T22444) / $signed(22'h100000);
  assign T22444 = $signed(31'h3fde0205) * $signed(16'hffff);
  assign T22445 = {T22448, T22446};
  assign T22446 = $signed(T22447) / $signed(22'h100000);
  assign T22447 = $signed(28'h41ed853) * $signed(16'h0);
  assign T22448 = T22449 ? 3'h7 : 3'h0;
  assign T22449 = T22446[6'h2b:6'h2b];
  assign T22450 = T18725[1'h0:1'h0];
  assign T22451 = T18725[1'h1:1'h1];
  assign T22452 = T22485 ? T22469 : T22453;
  assign T22453 = T22468 ? twiddle4_1_493_imag : twiddle4_1_492_imag;
  assign twiddle4_1_492_imag = T22456 + T22454;
  assign T22454 = $signed(T22455) / $signed(22'h100000);
  assign T22455 = $signed(31'h3fe12acb) * $signed(16'hffff);
  assign T22456 = {T22459, T22457};
  assign T22457 = $signed(T22458) / $signed(22'h100000);
  assign T22458 = $signed(27'h3ecadcf) * $signed(16'h0);
  assign T22459 = T22460 ? 4'hf : 4'h0;
  assign T22460 = T22457[6'h2a:6'h2a];
  assign twiddle4_1_493_imag = T22463 + T22461;
  assign T22461 = $signed(T22462) / $signed(22'h100000);
  assign T22462 = $signed(31'h3fe42c29) * $signed(16'hffff);
  assign T22463 = {T22466, T22464};
  assign T22464 = $signed(T22465) / $signed(22'h100000);
  assign T22465 = $signed(27'h3ba80df) * $signed(16'h0);
  assign T22466 = T22467 ? 4'hf : 4'h0;
  assign T22467 = T22464[6'h2a:6'h2a];
  assign T22468 = T18725[1'h0:1'h0];
  assign T22469 = T22484 ? twiddle4_1_495_imag : twiddle4_1_494_imag;
  assign twiddle4_1_494_imag = T22472 + T22470;
  assign T22470 = $signed(T22471) / $signed(22'h100000);
  assign T22471 = $signed(31'h3fe7061f) * $signed(16'hffff);
  assign T22472 = {T22475, T22473};
  assign T22473 = $signed(T22474) / $signed(22'h100000);
  assign T22474 = $signed(27'h38851a2) * $signed(16'h0);
  assign T22475 = T22476 ? 4'hf : 4'h0;
  assign T22476 = T22473[6'h2a:6'h2a];
  assign twiddle4_1_495_imag = T22479 + T22477;
  assign T22477 = $signed(T22478) / $signed(22'h100000);
  assign T22478 = $signed(31'h3fe9b8a9) * $signed(16'hffff);
  assign T22479 = {T22482, T22480};
  assign T22480 = $signed(T22481) / $signed(22'h100000);
  assign T22481 = $signed(27'h3562037) * $signed(16'h0);
  assign T22482 = T22483 ? 4'hf : 4'h0;
  assign T22483 = T22480[6'h2a:6'h2a];
  assign T22484 = T18725[1'h0:1'h0];
  assign T22485 = T18725[1'h1:1'h1];
  assign T22486 = T18725[2'h2:2'h2];
  assign T22487 = T18725[2'h3:2'h3];
  assign T22488 = T22629 ? T22559 : T22489;
  assign T22489 = T22558 ? T22524 : T22490;
  assign T22490 = T22523 ? T22507 : T22491;
  assign T22491 = T22506 ? twiddle4_1_497_imag : twiddle4_1_496_imag;
  assign twiddle4_1_496_imag = T22494 + T22492;
  assign T22492 = $signed(T22493) / $signed(22'h100000);
  assign T22493 = $signed(31'h3fec43c6) * $signed(16'hffff);
  assign T22494 = {T22497, T22495};
  assign T22495 = $signed(T22496) / $signed(22'h100000);
  assign T22496 = $signed(27'h323ecbe) * $signed(16'h0);
  assign T22497 = T22498 ? 4'hf : 4'h0;
  assign T22498 = T22495[6'h2a:6'h2a];
  assign twiddle4_1_497_imag = T22501 + T22499;
  assign T22499 = $signed(T22500) / $signed(22'h100000);
  assign T22500 = $signed(31'h3feea776) * $signed(16'hffff);
  assign T22501 = {T22504, T22502};
  assign T22502 = $signed(T22503) / $signed(22'h100000);
  assign T22503 = $signed(27'h2f1b754) * $signed(16'h0);
  assign T22504 = T22505 ? 4'hf : 4'h0;
  assign T22505 = T22502[6'h2a:6'h2a];
  assign T22506 = T18725[1'h0:1'h0];
  assign T22507 = T22522 ? twiddle4_1_499_imag : twiddle4_1_498_imag;
  assign twiddle4_1_498_imag = T22510 + T22508;
  assign T22508 = $signed(T22509) / $signed(22'h100000);
  assign T22509 = $signed(31'h3ff0e3b5) * $signed(16'hffff);
  assign T22510 = {T22513, T22511};
  assign T22511 = $signed(T22512) / $signed(22'h100000);
  assign T22512 = $signed(27'h2bf801a) * $signed(16'h0);
  assign T22513 = T22514 ? 4'hf : 4'h0;
  assign T22514 = T22511[6'h2a:6'h2a];
  assign twiddle4_1_499_imag = T22517 + T22515;
  assign T22515 = $signed(T22516) / $signed(22'h100000);
  assign T22516 = $signed(31'h3ff2f884) * $signed(16'hffff);
  assign T22517 = {T22520, T22518};
  assign T22518 = $signed(T22519) / $signed(22'h100000);
  assign T22519 = $signed(27'h28d472d) * $signed(16'h0);
  assign T22520 = T22521 ? 4'hf : 4'h0;
  assign T22521 = T22518[6'h2a:6'h2a];
  assign T22522 = T18725[1'h0:1'h0];
  assign T22523 = T18725[1'h1:1'h1];
  assign T22524 = T22557 ? T22541 : T22525;
  assign T22525 = T22540 ? twiddle4_1_501_imag : twiddle4_1_500_imag;
  assign twiddle4_1_500_imag = T22528 + T22526;
  assign T22526 = $signed(T22527) / $signed(22'h100000);
  assign T22527 = $signed(31'h3ff4e5df) * $signed(16'hffff);
  assign T22528 = {T22531, T22529};
  assign T22529 = $signed(T22530) / $signed(22'h100000);
  assign T22530 = $signed(27'h25b0cae) * $signed(16'h0);
  assign T22531 = T22532 ? 4'hf : 4'h0;
  assign T22532 = T22529[6'h2a:6'h2a];
  assign twiddle4_1_501_imag = T22535 + T22533;
  assign T22533 = $signed(T22534) / $signed(22'h100000);
  assign T22534 = $signed(31'h3ff6abc8) * $signed(16'hffff);
  assign T22535 = {T22538, T22536};
  assign T22536 = $signed(T22537) / $signed(22'h100000);
  assign T22537 = $signed(27'h228d0bb) * $signed(16'h0);
  assign T22538 = T22539 ? 4'hf : 4'h0;
  assign T22539 = T22536[6'h2a:6'h2a];
  assign T22540 = T18725[1'h0:1'h0];
  assign T22541 = T22556 ? twiddle4_1_503_imag : twiddle4_1_502_imag;
  assign twiddle4_1_502_imag = T22544 + T22542;
  assign T22542 = $signed(T22543) / $signed(22'h100000);
  assign T22543 = $signed(31'h3ff84a3b) * $signed(16'hffff);
  assign T22544 = {T22547, T22545};
  assign T22545 = $signed(T22546) / $signed(22'h100000);
  assign T22546 = $signed(26'h1f69373) * $signed(16'h0);
  assign T22547 = T22548 ? 5'h1f : 5'h0;
  assign T22548 = T22545[6'h29:6'h29];
  assign twiddle4_1_503_imag = T22551 + T22549;
  assign T22549 = $signed(T22550) / $signed(22'h100000);
  assign T22550 = $signed(31'h3ff9c139) * $signed(16'hffff);
  assign T22551 = {T22554, T22552};
  assign T22552 = $signed(T22553) / $signed(22'h100000);
  assign T22553 = $signed(26'h1c454f4) * $signed(16'h0);
  assign T22554 = T22555 ? 5'h1f : 5'h0;
  assign T22555 = T22552[6'h29:6'h29];
  assign T22556 = T18725[1'h0:1'h0];
  assign T22557 = T18725[1'h1:1'h1];
  assign T22558 = T18725[2'h2:2'h2];
  assign T22559 = T22628 ? T22594 : T22560;
  assign T22560 = T22593 ? T22577 : T22561;
  assign T22561 = T22576 ? twiddle4_1_505_imag : twiddle4_1_504_imag;
  assign twiddle4_1_504_imag = T22564 + T22562;
  assign T22562 = $signed(T22563) / $signed(22'h100000);
  assign T22563 = $signed(31'h3ffb10c1) * $signed(16'hffff);
  assign T22564 = {T22567, T22565};
  assign T22565 = $signed(T22566) / $signed(22'h100000);
  assign T22566 = $signed(26'h192155f) * $signed(16'h0);
  assign T22567 = T22568 ? 5'h1f : 5'h0;
  assign T22568 = T22565[6'h29:6'h29];
  assign twiddle4_1_505_imag = T22571 + T22569;
  assign T22569 = $signed(T22570) / $signed(22'h100000);
  assign T22570 = $signed(31'h3ffc38d0) * $signed(16'hffff);
  assign T22571 = {T22574, T22572};
  assign T22572 = $signed(T22573) / $signed(22'h100000);
  assign T22573 = $signed(26'h15fd4d2) * $signed(16'h0);
  assign T22574 = T22575 ? 5'h1f : 5'h0;
  assign T22575 = T22572[6'h29:6'h29];
  assign T22576 = T18725[1'h0:1'h0];
  assign T22577 = T22592 ? twiddle4_1_507_imag : twiddle4_1_506_imag;
  assign twiddle4_1_506_imag = T22580 + T22578;
  assign T22578 = $signed(T22579) / $signed(22'h100000);
  assign T22579 = $signed(31'h3ffd3968) * $signed(16'hffff);
  assign T22580 = {T22583, T22581};
  assign T22581 = $signed(T22582) / $signed(22'h100000);
  assign T22582 = $signed(26'h12d936b) * $signed(16'h0);
  assign T22583 = T22584 ? 5'h1f : 5'h0;
  assign T22584 = T22581[6'h29:6'h29];
  assign twiddle4_1_507_imag = T22587 + T22585;
  assign T22585 = $signed(T22586) / $signed(22'h100000);
  assign T22586 = $signed(31'h3ffe1287) * $signed(16'hffff);
  assign T22587 = {T22590, T22588};
  assign T22588 = $signed(T22589) / $signed(22'h100000);
  assign T22589 = $signed(25'hfb514b) * $signed(16'h0);
  assign T22590 = T22591 ? 6'h3f : 6'h0;
  assign T22591 = T22588[6'h28:6'h28];
  assign T22592 = T18725[1'h0:1'h0];
  assign T22593 = T18725[1'h1:1'h1];
  assign T22594 = T22627 ? T22611 : T22595;
  assign T22595 = T22610 ? twiddle4_1_509_imag : twiddle4_1_508_imag;
  assign twiddle4_1_508_imag = T22598 + T22596;
  assign T22596 = $signed(T22597) / $signed(22'h100000);
  assign T22597 = $signed(31'h3ffec42d) * $signed(16'hffff);
  assign T22598 = {T22601, T22599};
  assign T22599 = $signed(T22600) / $signed(22'h100000);
  assign T22600 = $signed(25'hc90e8f) * $signed(16'h0);
  assign T22601 = T22602 ? 6'h3f : 6'h0;
  assign T22602 = T22599[6'h28:6'h28];
  assign twiddle4_1_509_imag = T22605 + T22603;
  assign T22603 = $signed(T22604) / $signed(22'h100000);
  assign T22604 = $signed(31'h3fff4e59) * $signed(16'hffff);
  assign T22605 = {T22608, T22606};
  assign T22606 = $signed(T22607) / $signed(22'h100000);
  assign T22607 = $signed(25'h96cb58) * $signed(16'h0);
  assign T22608 = T22609 ? 6'h3f : 6'h0;
  assign T22609 = T22606[6'h28:6'h28];
  assign T22610 = T18725[1'h0:1'h0];
  assign T22611 = T22626 ? twiddle4_1_511_imag : twiddle4_1_510_imag;
  assign twiddle4_1_510_imag = T22614 + T22612;
  assign T22612 = $signed(T22613) / $signed(22'h100000);
  assign T22613 = $signed(31'h3fffb10b) * $signed(16'hffff);
  assign T22614 = {T22617, T22615};
  assign T22615 = $signed(T22616) / $signed(22'h100000);
  assign T22616 = $signed(24'h6487c3) * $signed(16'h0);
  assign T22617 = T22618 ? 7'h7f : 7'h0;
  assign T22618 = T22615[6'h27:6'h27];
  assign twiddle4_1_511_imag = T22621 + T22619;
  assign T22619 = $signed(T22620) / $signed(22'h100000);
  assign T22620 = $signed(31'h3fffec42) * $signed(16'hffff);
  assign T22621 = {T22624, T22622};
  assign T22622 = $signed(T22623) / $signed(22'h100000);
  assign T22623 = $signed(23'h3243f1) * $signed(16'h0);
  assign T22624 = T22625 ? 8'hff : 8'h0;
  assign T22625 = T22622[6'h26:6'h26];
  assign T22626 = T18725[1'h0:1'h0];
  assign T22627 = T18725[1'h1:1'h1];
  assign T22628 = T18725[2'h2:2'h2];
  assign T22629 = T18725[2'h3:2'h3];
  assign T22630 = T18725[3'h4:3'h4];
  assign T22631 = T18725[3'h5:3'h5];
  assign T22632 = T18725[3'h6:3'h6];
  assign T22633 = T18725[3'h7:3'h7];
  assign T22634 = T20678[6'h2e:6'h2e];
  assign T22635 = T18725[4'h8:4'h8];
  assign io_t4_1out_real = T22636;
  assign T22636 = T22637[4'hf:1'h0];
  assign T22637 = T26571 ? T24613 : T22638;
  assign T22638 = T24612 ? T23758 : T22639;
  assign T22639 = T23757 ? T23226 : T22640;
  assign T22640 = T23225 ? T22937 : T22641;
  assign T22641 = T22936 ? T22792 : T22642;
  assign T22642 = T22791 ? T22719 : T22643;
  assign T22643 = T22718 ? T22682 : T22644;
  assign T22644 = T22681 ? T22663 : T22645;
  assign T22645 = T22662 ? T22653 : twiddle4_1_0_real;
  assign twiddle4_1_0_real = T22651 + T22646;
  assign T22646 = {T22649, T22647};
  assign T22647 = $signed(T22648) / $signed(22'h100000);
  assign T22648 = $signed(1'h0) * $signed(16'h0);
  assign T22649 = T22650 ? 31'h7fffffff : 31'h0;
  assign T22650 = T22647[5'h10:5'h10];
  assign T22651 = $signed(T22652) / $signed(22'h100000);
  assign T22652 = $signed(32'h40000000) * $signed(16'h1);
  assign T22653 = {T22661, twiddle4_1_1_real};
  assign twiddle4_1_1_real = T22659 + T22654;
  assign T22654 = {T22657, T22655};
  assign T22655 = $signed(T22656) / $signed(22'h100000);
  assign T22656 = $signed(23'h3243f1) * $signed(16'h0);
  assign T22657 = T22658 ? 8'hff : 8'h0;
  assign T22658 = T22655[6'h26:6'h26];
  assign T22659 = $signed(T22660) / $signed(22'h100000);
  assign T22660 = $signed(31'h3fffec42) * $signed(16'h1);
  assign T22661 = twiddle4_1_1_real[6'h2e:6'h2e];
  assign T22662 = T18725[1'h0:1'h0];
  assign T22663 = {T22680, T22664};
  assign T22664 = T22679 ? twiddle4_1_3_real : twiddle4_1_2_real;
  assign twiddle4_1_2_real = T22670 + T22665;
  assign T22665 = {T22668, T22666};
  assign T22666 = $signed(T22667) / $signed(22'h100000);
  assign T22667 = $signed(24'h6487c3) * $signed(16'h0);
  assign T22668 = T22669 ? 7'h7f : 7'h0;
  assign T22669 = T22666[6'h27:6'h27];
  assign T22670 = $signed(T22671) / $signed(22'h100000);
  assign T22671 = $signed(31'h3fffb10b) * $signed(16'h1);
  assign twiddle4_1_3_real = T22677 + T22672;
  assign T22672 = {T22675, T22673};
  assign T22673 = $signed(T22674) / $signed(22'h100000);
  assign T22674 = $signed(25'h96cb58) * $signed(16'h0);
  assign T22675 = T22676 ? 6'h3f : 6'h0;
  assign T22676 = T22673[6'h28:6'h28];
  assign T22677 = $signed(T22678) / $signed(22'h100000);
  assign T22678 = $signed(31'h3fff4e59) * $signed(16'h1);
  assign T22679 = T18725[1'h0:1'h0];
  assign T22680 = T22664[6'h2e:6'h2e];
  assign T22681 = T18725[1'h1:1'h1];
  assign T22682 = {T22717, T22683};
  assign T22683 = T22716 ? T22700 : T22684;
  assign T22684 = T22699 ? twiddle4_1_5_real : twiddle4_1_4_real;
  assign twiddle4_1_4_real = T22690 + T22685;
  assign T22685 = {T22688, T22686};
  assign T22686 = $signed(T22687) / $signed(22'h100000);
  assign T22687 = $signed(25'hc90e8f) * $signed(16'h0);
  assign T22688 = T22689 ? 6'h3f : 6'h0;
  assign T22689 = T22686[6'h28:6'h28];
  assign T22690 = $signed(T22691) / $signed(22'h100000);
  assign T22691 = $signed(31'h3ffec42d) * $signed(16'h1);
  assign twiddle4_1_5_real = T22697 + T22692;
  assign T22692 = {T22695, T22693};
  assign T22693 = $signed(T22694) / $signed(22'h100000);
  assign T22694 = $signed(25'hfb514b) * $signed(16'h0);
  assign T22695 = T22696 ? 6'h3f : 6'h0;
  assign T22696 = T22693[6'h28:6'h28];
  assign T22697 = $signed(T22698) / $signed(22'h100000);
  assign T22698 = $signed(31'h3ffe1287) * $signed(16'h1);
  assign T22699 = T18725[1'h0:1'h0];
  assign T22700 = T22715 ? twiddle4_1_7_real : twiddle4_1_6_real;
  assign twiddle4_1_6_real = T22706 + T22701;
  assign T22701 = {T22704, T22702};
  assign T22702 = $signed(T22703) / $signed(22'h100000);
  assign T22703 = $signed(26'h12d936b) * $signed(16'h0);
  assign T22704 = T22705 ? 5'h1f : 5'h0;
  assign T22705 = T22702[6'h29:6'h29];
  assign T22706 = $signed(T22707) / $signed(22'h100000);
  assign T22707 = $signed(31'h3ffd3968) * $signed(16'h1);
  assign twiddle4_1_7_real = T22713 + T22708;
  assign T22708 = {T22711, T22709};
  assign T22709 = $signed(T22710) / $signed(22'h100000);
  assign T22710 = $signed(26'h15fd4d2) * $signed(16'h0);
  assign T22711 = T22712 ? 5'h1f : 5'h0;
  assign T22712 = T22709[6'h29:6'h29];
  assign T22713 = $signed(T22714) / $signed(22'h100000);
  assign T22714 = $signed(31'h3ffc38d0) * $signed(16'h1);
  assign T22715 = T18725[1'h0:1'h0];
  assign T22716 = T18725[1'h1:1'h1];
  assign T22717 = T22683[6'h2e:6'h2e];
  assign T22718 = T18725[2'h2:2'h2];
  assign T22719 = {T22790, T22720};
  assign T22720 = T22789 ? T22755 : T22721;
  assign T22721 = T22754 ? T22738 : T22722;
  assign T22722 = T22737 ? twiddle4_1_9_real : twiddle4_1_8_real;
  assign twiddle4_1_8_real = T22728 + T22723;
  assign T22723 = {T22726, T22724};
  assign T22724 = $signed(T22725) / $signed(22'h100000);
  assign T22725 = $signed(26'h192155f) * $signed(16'h0);
  assign T22726 = T22727 ? 5'h1f : 5'h0;
  assign T22727 = T22724[6'h29:6'h29];
  assign T22728 = $signed(T22729) / $signed(22'h100000);
  assign T22729 = $signed(31'h3ffb10c1) * $signed(16'h1);
  assign twiddle4_1_9_real = T22735 + T22730;
  assign T22730 = {T22733, T22731};
  assign T22731 = $signed(T22732) / $signed(22'h100000);
  assign T22732 = $signed(26'h1c454f4) * $signed(16'h0);
  assign T22733 = T22734 ? 5'h1f : 5'h0;
  assign T22734 = T22731[6'h29:6'h29];
  assign T22735 = $signed(T22736) / $signed(22'h100000);
  assign T22736 = $signed(31'h3ff9c139) * $signed(16'h1);
  assign T22737 = T18725[1'h0:1'h0];
  assign T22738 = T22753 ? twiddle4_1_11_real : twiddle4_1_10_real;
  assign twiddle4_1_10_real = T22744 + T22739;
  assign T22739 = {T22742, T22740};
  assign T22740 = $signed(T22741) / $signed(22'h100000);
  assign T22741 = $signed(26'h1f69373) * $signed(16'h0);
  assign T22742 = T22743 ? 5'h1f : 5'h0;
  assign T22743 = T22740[6'h29:6'h29];
  assign T22744 = $signed(T22745) / $signed(22'h100000);
  assign T22745 = $signed(31'h3ff84a3b) * $signed(16'h1);
  assign twiddle4_1_11_real = T22751 + T22746;
  assign T22746 = {T22749, T22747};
  assign T22747 = $signed(T22748) / $signed(22'h100000);
  assign T22748 = $signed(27'h228d0bb) * $signed(16'h0);
  assign T22749 = T22750 ? 4'hf : 4'h0;
  assign T22750 = T22747[6'h2a:6'h2a];
  assign T22751 = $signed(T22752) / $signed(22'h100000);
  assign T22752 = $signed(31'h3ff6abc8) * $signed(16'h1);
  assign T22753 = T18725[1'h0:1'h0];
  assign T22754 = T18725[1'h1:1'h1];
  assign T22755 = T22788 ? T22772 : T22756;
  assign T22756 = T22771 ? twiddle4_1_13_real : twiddle4_1_12_real;
  assign twiddle4_1_12_real = T22762 + T22757;
  assign T22757 = {T22760, T22758};
  assign T22758 = $signed(T22759) / $signed(22'h100000);
  assign T22759 = $signed(27'h25b0cae) * $signed(16'h0);
  assign T22760 = T22761 ? 4'hf : 4'h0;
  assign T22761 = T22758[6'h2a:6'h2a];
  assign T22762 = $signed(T22763) / $signed(22'h100000);
  assign T22763 = $signed(31'h3ff4e5df) * $signed(16'h1);
  assign twiddle4_1_13_real = T22769 + T22764;
  assign T22764 = {T22767, T22765};
  assign T22765 = $signed(T22766) / $signed(22'h100000);
  assign T22766 = $signed(27'h28d472d) * $signed(16'h0);
  assign T22767 = T22768 ? 4'hf : 4'h0;
  assign T22768 = T22765[6'h2a:6'h2a];
  assign T22769 = $signed(T22770) / $signed(22'h100000);
  assign T22770 = $signed(31'h3ff2f884) * $signed(16'h1);
  assign T22771 = T18725[1'h0:1'h0];
  assign T22772 = T22787 ? twiddle4_1_15_real : twiddle4_1_14_real;
  assign twiddle4_1_14_real = T22778 + T22773;
  assign T22773 = {T22776, T22774};
  assign T22774 = $signed(T22775) / $signed(22'h100000);
  assign T22775 = $signed(27'h2bf801a) * $signed(16'h0);
  assign T22776 = T22777 ? 4'hf : 4'h0;
  assign T22777 = T22774[6'h2a:6'h2a];
  assign T22778 = $signed(T22779) / $signed(22'h100000);
  assign T22779 = $signed(31'h3ff0e3b5) * $signed(16'h1);
  assign twiddle4_1_15_real = T22785 + T22780;
  assign T22780 = {T22783, T22781};
  assign T22781 = $signed(T22782) / $signed(22'h100000);
  assign T22782 = $signed(27'h2f1b754) * $signed(16'h0);
  assign T22783 = T22784 ? 4'hf : 4'h0;
  assign T22784 = T22781[6'h2a:6'h2a];
  assign T22785 = $signed(T22786) / $signed(22'h100000);
  assign T22786 = $signed(31'h3feea776) * $signed(16'h1);
  assign T22787 = T18725[1'h0:1'h0];
  assign T22788 = T18725[1'h1:1'h1];
  assign T22789 = T18725[2'h2:2'h2];
  assign T22790 = T22720[6'h2e:6'h2e];
  assign T22791 = T18725[2'h3:2'h3];
  assign T22792 = {T22935, T22793};
  assign T22793 = T22934 ? T22864 : T22794;
  assign T22794 = T22863 ? T22829 : T22795;
  assign T22795 = T22828 ? T22812 : T22796;
  assign T22796 = T22811 ? twiddle4_1_17_real : twiddle4_1_16_real;
  assign twiddle4_1_16_real = T22802 + T22797;
  assign T22797 = {T22800, T22798};
  assign T22798 = $signed(T22799) / $signed(22'h100000);
  assign T22799 = $signed(27'h323ecbe) * $signed(16'h0);
  assign T22800 = T22801 ? 4'hf : 4'h0;
  assign T22801 = T22798[6'h2a:6'h2a];
  assign T22802 = $signed(T22803) / $signed(22'h100000);
  assign T22803 = $signed(31'h3fec43c6) * $signed(16'h1);
  assign twiddle4_1_17_real = T22809 + T22804;
  assign T22804 = {T22807, T22805};
  assign T22805 = $signed(T22806) / $signed(22'h100000);
  assign T22806 = $signed(27'h3562037) * $signed(16'h0);
  assign T22807 = T22808 ? 4'hf : 4'h0;
  assign T22808 = T22805[6'h2a:6'h2a];
  assign T22809 = $signed(T22810) / $signed(22'h100000);
  assign T22810 = $signed(31'h3fe9b8a9) * $signed(16'h1);
  assign T22811 = T18725[1'h0:1'h0];
  assign T22812 = T22827 ? twiddle4_1_19_real : twiddle4_1_18_real;
  assign twiddle4_1_18_real = T22818 + T22813;
  assign T22813 = {T22816, T22814};
  assign T22814 = $signed(T22815) / $signed(22'h100000);
  assign T22815 = $signed(27'h38851a2) * $signed(16'h0);
  assign T22816 = T22817 ? 4'hf : 4'h0;
  assign T22817 = T22814[6'h2a:6'h2a];
  assign T22818 = $signed(T22819) / $signed(22'h100000);
  assign T22819 = $signed(31'h3fe7061f) * $signed(16'h1);
  assign twiddle4_1_19_real = T22825 + T22820;
  assign T22820 = {T22823, T22821};
  assign T22821 = $signed(T22822) / $signed(22'h100000);
  assign T22822 = $signed(27'h3ba80df) * $signed(16'h0);
  assign T22823 = T22824 ? 4'hf : 4'h0;
  assign T22824 = T22821[6'h2a:6'h2a];
  assign T22825 = $signed(T22826) / $signed(22'h100000);
  assign T22826 = $signed(31'h3fe42c29) * $signed(16'h1);
  assign T22827 = T18725[1'h0:1'h0];
  assign T22828 = T18725[1'h1:1'h1];
  assign T22829 = T22862 ? T22846 : T22830;
  assign T22830 = T22845 ? twiddle4_1_21_real : twiddle4_1_20_real;
  assign twiddle4_1_20_real = T22836 + T22831;
  assign T22831 = {T22834, T22832};
  assign T22832 = $signed(T22833) / $signed(22'h100000);
  assign T22833 = $signed(27'h3ecadcf) * $signed(16'h0);
  assign T22834 = T22835 ? 4'hf : 4'h0;
  assign T22835 = T22832[6'h2a:6'h2a];
  assign T22836 = $signed(T22837) / $signed(22'h100000);
  assign T22837 = $signed(31'h3fe12acb) * $signed(16'h1);
  assign twiddle4_1_21_real = T22843 + T22838;
  assign T22838 = {T22841, T22839};
  assign T22839 = $signed(T22840) / $signed(22'h100000);
  assign T22840 = $signed(28'h41ed853) * $signed(16'h0);
  assign T22841 = T22842 ? 3'h7 : 3'h0;
  assign T22842 = T22839[6'h2b:6'h2b];
  assign T22843 = $signed(T22844) / $signed(22'h100000);
  assign T22844 = $signed(31'h3fde0205) * $signed(16'h1);
  assign T22845 = T18725[1'h0:1'h0];
  assign T22846 = T22861 ? twiddle4_1_23_real : twiddle4_1_22_real;
  assign twiddle4_1_22_real = T22852 + T22847;
  assign T22847 = {T22850, T22848};
  assign T22848 = $signed(T22849) / $signed(22'h100000);
  assign T22849 = $signed(28'h451004d) * $signed(16'h0);
  assign T22850 = T22851 ? 3'h7 : 3'h0;
  assign T22851 = T22848[6'h2b:6'h2b];
  assign T22852 = $signed(T22853) / $signed(22'h100000);
  assign T22853 = $signed(31'h3fdab1d9) * $signed(16'h1);
  assign twiddle4_1_23_real = T22859 + T22854;
  assign T22854 = {T22857, T22855};
  assign T22855 = $signed(T22856) / $signed(22'h100000);
  assign T22856 = $signed(28'h483259d) * $signed(16'h0);
  assign T22857 = T22858 ? 3'h7 : 3'h0;
  assign T22858 = T22855[6'h2b:6'h2b];
  assign T22859 = $signed(T22860) / $signed(22'h100000);
  assign T22860 = $signed(31'h3fd73a4a) * $signed(16'h1);
  assign T22861 = T18725[1'h0:1'h0];
  assign T22862 = T18725[1'h1:1'h1];
  assign T22863 = T18725[2'h2:2'h2];
  assign T22864 = T22933 ? T22899 : T22865;
  assign T22865 = T22898 ? T22882 : T22866;
  assign T22866 = T22881 ? twiddle4_1_25_real : twiddle4_1_24_real;
  assign twiddle4_1_24_real = T22872 + T22867;
  assign T22867 = {T22870, T22868};
  assign T22868 = $signed(T22869) / $signed(22'h100000);
  assign T22869 = $signed(28'h4b54824) * $signed(16'h0);
  assign T22870 = T22871 ? 3'h7 : 3'h0;
  assign T22871 = T22868[6'h2b:6'h2b];
  assign T22872 = $signed(T22873) / $signed(22'h100000);
  assign T22873 = $signed(31'h3fd39b5a) * $signed(16'h1);
  assign twiddle4_1_25_real = T22879 + T22874;
  assign T22874 = {T22877, T22875};
  assign T22875 = $signed(T22876) / $signed(22'h100000);
  assign T22876 = $signed(28'h4e767c4) * $signed(16'h0);
  assign T22877 = T22878 ? 3'h7 : 3'h0;
  assign T22878 = T22875[6'h2b:6'h2b];
  assign T22879 = $signed(T22880) / $signed(22'h100000);
  assign T22880 = $signed(31'h3fcfd50a) * $signed(16'h1);
  assign T22881 = T18725[1'h0:1'h0];
  assign T22882 = T22897 ? twiddle4_1_27_real : twiddle4_1_26_real;
  assign twiddle4_1_26_real = T22888 + T22883;
  assign T22883 = {T22886, T22884};
  assign T22884 = $signed(T22885) / $signed(22'h100000);
  assign T22885 = $signed(28'h519845e) * $signed(16'h0);
  assign T22886 = T22887 ? 3'h7 : 3'h0;
  assign T22887 = T22884[6'h2b:6'h2b];
  assign T22888 = $signed(T22889) / $signed(22'h100000);
  assign T22889 = $signed(31'h3fcbe75e) * $signed(16'h1);
  assign twiddle4_1_27_real = T22895 + T22890;
  assign T22890 = {T22893, T22891};
  assign T22891 = $signed(T22892) / $signed(22'h100000);
  assign T22892 = $signed(28'h54b9dd2) * $signed(16'h0);
  assign T22893 = T22894 ? 3'h7 : 3'h0;
  assign T22894 = T22891[6'h2b:6'h2b];
  assign T22895 = $signed(T22896) / $signed(22'h100000);
  assign T22896 = $signed(31'h3fc7d257) * $signed(16'h1);
  assign T22897 = T18725[1'h0:1'h0];
  assign T22898 = T18725[1'h1:1'h1];
  assign T22899 = T22932 ? T22916 : T22900;
  assign T22900 = T22915 ? twiddle4_1_29_real : twiddle4_1_28_real;
  assign twiddle4_1_28_real = T22906 + T22901;
  assign T22901 = {T22904, T22902};
  assign T22902 = $signed(T22903) / $signed(22'h100000);
  assign T22903 = $signed(28'h57db402) * $signed(16'h0);
  assign T22904 = T22905 ? 3'h7 : 3'h0;
  assign T22905 = T22902[6'h2b:6'h2b];
  assign T22906 = $signed(T22907) / $signed(22'h100000);
  assign T22907 = $signed(31'h3fc395f9) * $signed(16'h1);
  assign twiddle4_1_29_real = T22913 + T22908;
  assign T22908 = {T22911, T22909};
  assign T22909 = $signed(T22910) / $signed(22'h100000);
  assign T22910 = $signed(28'h5afc6cf) * $signed(16'h0);
  assign T22911 = T22912 ? 3'h7 : 3'h0;
  assign T22912 = T22909[6'h2b:6'h2b];
  assign T22913 = $signed(T22914) / $signed(22'h100000);
  assign T22914 = $signed(31'h3fbf3245) * $signed(16'h1);
  assign T22915 = T18725[1'h0:1'h0];
  assign T22916 = T22931 ? twiddle4_1_31_real : twiddle4_1_30_real;
  assign twiddle4_1_30_real = T22922 + T22917;
  assign T22917 = {T22920, T22918};
  assign T22918 = $signed(T22919) / $signed(22'h100000);
  assign T22919 = $signed(28'h5e1d61a) * $signed(16'h0);
  assign T22920 = T22921 ? 3'h7 : 3'h0;
  assign T22921 = T22918[6'h2b:6'h2b];
  assign T22922 = $signed(T22923) / $signed(22'h100000);
  assign T22923 = $signed(31'h3fbaa73f) * $signed(16'h1);
  assign twiddle4_1_31_real = T22929 + T22924;
  assign T22924 = {T22927, T22925};
  assign T22925 = $signed(T22926) / $signed(22'h100000);
  assign T22926 = $signed(28'h613e1c4) * $signed(16'h0);
  assign T22927 = T22928 ? 3'h7 : 3'h0;
  assign T22928 = T22925[6'h2b:6'h2b];
  assign T22929 = $signed(T22930) / $signed(22'h100000);
  assign T22930 = $signed(31'h3fb5f4ea) * $signed(16'h1);
  assign T22931 = T18725[1'h0:1'h0];
  assign T22932 = T18725[1'h1:1'h1];
  assign T22933 = T18725[2'h2:2'h2];
  assign T22934 = T18725[2'h3:2'h3];
  assign T22935 = T22793[6'h2e:6'h2e];
  assign T22936 = T18725[3'h4:3'h4];
  assign T22937 = {T23224, T22938};
  assign T22938 = T23223 ? T23081 : T22939;
  assign T22939 = T23080 ? T23010 : T22940;
  assign T22940 = T23009 ? T22975 : T22941;
  assign T22941 = T22974 ? T22958 : T22942;
  assign T22942 = T22957 ? twiddle4_1_33_real : twiddle4_1_32_real;
  assign twiddle4_1_32_real = T22948 + T22943;
  assign T22943 = {T22946, T22944};
  assign T22944 = $signed(T22945) / $signed(22'h100000);
  assign T22945 = $signed(28'h645e9af) * $signed(16'h0);
  assign T22946 = T22947 ? 3'h7 : 3'h0;
  assign T22947 = T22944[6'h2b:6'h2b];
  assign T22948 = $signed(T22949) / $signed(22'h100000);
  assign T22949 = $signed(31'h3fb11b47) * $signed(16'h1);
  assign twiddle4_1_33_real = T22955 + T22950;
  assign T22950 = {T22953, T22951};
  assign T22951 = $signed(T22952) / $signed(22'h100000);
  assign T22952 = $signed(28'h677edba) * $signed(16'h0);
  assign T22953 = T22954 ? 3'h7 : 3'h0;
  assign T22954 = T22951[6'h2b:6'h2b];
  assign T22955 = $signed(T22956) / $signed(22'h100000);
  assign T22956 = $signed(31'h3fac1a5b) * $signed(16'h1);
  assign T22957 = T18725[1'h0:1'h0];
  assign T22958 = T22973 ? twiddle4_1_35_real : twiddle4_1_34_real;
  assign twiddle4_1_34_real = T22964 + T22959;
  assign T22959 = {T22962, T22960};
  assign T22960 = $signed(T22961) / $signed(22'h100000);
  assign T22961 = $signed(28'h6a9edc9) * $signed(16'h0);
  assign T22962 = T22963 ? 3'h7 : 3'h0;
  assign T22963 = T22960[6'h2b:6'h2b];
  assign T22964 = $signed(T22965) / $signed(22'h100000);
  assign T22965 = $signed(31'h3fa6f228) * $signed(16'h1);
  assign twiddle4_1_35_real = T22971 + T22966;
  assign T22966 = {T22969, T22967};
  assign T22967 = $signed(T22968) / $signed(22'h100000);
  assign T22968 = $signed(28'h6dbe9bb) * $signed(16'h0);
  assign T22969 = T22970 ? 3'h7 : 3'h0;
  assign T22970 = T22967[6'h2b:6'h2b];
  assign T22971 = $signed(T22972) / $signed(22'h100000);
  assign T22972 = $signed(31'h3fa1a2b1) * $signed(16'h1);
  assign T22973 = T18725[1'h0:1'h0];
  assign T22974 = T18725[1'h1:1'h1];
  assign T22975 = T23008 ? T22992 : T22976;
  assign T22976 = T22991 ? twiddle4_1_37_real : twiddle4_1_36_real;
  assign twiddle4_1_36_real = T22982 + T22977;
  assign T22977 = {T22980, T22978};
  assign T22978 = $signed(T22979) / $signed(22'h100000);
  assign T22979 = $signed(28'h70de171) * $signed(16'h0);
  assign T22980 = T22981 ? 3'h7 : 3'h0;
  assign T22981 = T22978[6'h2b:6'h2b];
  assign T22982 = $signed(T22983) / $signed(22'h100000);
  assign T22983 = $signed(31'h3f9c2bfa) * $signed(16'h1);
  assign twiddle4_1_37_real = T22989 + T22984;
  assign T22984 = {T22987, T22985};
  assign T22985 = $signed(T22986) / $signed(22'h100000);
  assign T22986 = $signed(28'h73fd4ce) * $signed(16'h0);
  assign T22987 = T22988 ? 3'h7 : 3'h0;
  assign T22988 = T22985[6'h2b:6'h2b];
  assign T22989 = $signed(T22990) / $signed(22'h100000);
  assign T22990 = $signed(31'h3f968e07) * $signed(16'h1);
  assign T22991 = T18725[1'h0:1'h0];
  assign T22992 = T23007 ? twiddle4_1_39_real : twiddle4_1_38_real;
  assign twiddle4_1_38_real = T22998 + T22993;
  assign T22993 = {T22996, T22994};
  assign T22994 = $signed(T22995) / $signed(22'h100000);
  assign T22995 = $signed(28'h771c3b2) * $signed(16'h0);
  assign T22996 = T22997 ? 3'h7 : 3'h0;
  assign T22997 = T22994[6'h2b:6'h2b];
  assign T22998 = $signed(T22999) / $signed(22'h100000);
  assign T22999 = $signed(31'h3f90c8d9) * $signed(16'h1);
  assign twiddle4_1_39_real = T23005 + T23000;
  assign T23000 = {T23003, T23001};
  assign T23001 = $signed(T23002) / $signed(22'h100000);
  assign T23002 = $signed(28'h7a3adff) * $signed(16'h0);
  assign T23003 = T23004 ? 3'h7 : 3'h0;
  assign T23004 = T23001[6'h2b:6'h2b];
  assign T23005 = $signed(T23006) / $signed(22'h100000);
  assign T23006 = $signed(31'h3f8adc76) * $signed(16'h1);
  assign T23007 = T18725[1'h0:1'h0];
  assign T23008 = T18725[1'h1:1'h1];
  assign T23009 = T18725[2'h2:2'h2];
  assign T23010 = T23079 ? T23045 : T23011;
  assign T23011 = T23044 ? T23028 : T23012;
  assign T23012 = T23027 ? twiddle4_1_41_real : twiddle4_1_40_real;
  assign twiddle4_1_40_real = T23018 + T23013;
  assign T23013 = {T23016, T23014};
  assign T23014 = $signed(T23015) / $signed(22'h100000);
  assign T23015 = $signed(28'h7d59395) * $signed(16'h0);
  assign T23016 = T23017 ? 3'h7 : 3'h0;
  assign T23017 = T23014[6'h2b:6'h2b];
  assign T23018 = $signed(T23019) / $signed(22'h100000);
  assign T23019 = $signed(31'h3f84c8e1) * $signed(16'h1);
  assign twiddle4_1_41_real = T23025 + T23020;
  assign T23020 = {T23023, T23021};
  assign T23021 = $signed(T23022) / $signed(22'h100000);
  assign T23022 = $signed(29'h8077456) * $signed(16'h0);
  assign T23023 = T23024 ? 2'h3 : 2'h0;
  assign T23024 = T23021[6'h2c:6'h2c];
  assign T23025 = $signed(T23026) / $signed(22'h100000);
  assign T23026 = $signed(31'h3f7e8e1e) * $signed(16'h1);
  assign T23027 = T18725[1'h0:1'h0];
  assign T23028 = T23043 ? twiddle4_1_43_real : twiddle4_1_42_real;
  assign twiddle4_1_42_real = T23034 + T23029;
  assign T23029 = {T23032, T23030};
  assign T23030 = $signed(T23031) / $signed(22'h100000);
  assign T23031 = $signed(29'h8395023) * $signed(16'h0);
  assign T23032 = T23033 ? 2'h3 : 2'h0;
  assign T23033 = T23030[6'h2c:6'h2c];
  assign T23034 = $signed(T23035) / $signed(22'h100000);
  assign T23035 = $signed(31'h3f782c2f) * $signed(16'h1);
  assign twiddle4_1_43_real = T23041 + T23036;
  assign T23036 = {T23039, T23037};
  assign T23037 = $signed(T23038) / $signed(22'h100000);
  assign T23038 = $signed(29'h86b26de) * $signed(16'h0);
  assign T23039 = T23040 ? 2'h3 : 2'h0;
  assign T23040 = T23037[6'h2c:6'h2c];
  assign T23041 = $signed(T23042) / $signed(22'h100000);
  assign T23042 = $signed(31'h3f71a31a) * $signed(16'h1);
  assign T23043 = T18725[1'h0:1'h0];
  assign T23044 = T18725[1'h1:1'h1];
  assign T23045 = T23078 ? T23062 : T23046;
  assign T23046 = T23061 ? twiddle4_1_45_real : twiddle4_1_44_real;
  assign twiddle4_1_44_real = T23052 + T23047;
  assign T23047 = {T23050, T23048};
  assign T23048 = $signed(T23049) / $signed(22'h100000);
  assign T23049 = $signed(29'h89cf867) * $signed(16'h0);
  assign T23050 = T23051 ? 2'h3 : 2'h0;
  assign T23051 = T23048[6'h2c:6'h2c];
  assign T23052 = $signed(T23053) / $signed(22'h100000);
  assign T23053 = $signed(31'h3f6af2e3) * $signed(16'h1);
  assign twiddle4_1_45_real = T23059 + T23054;
  assign T23054 = {T23057, T23055};
  assign T23055 = $signed(T23056) / $signed(22'h100000);
  assign T23056 = $signed(29'h8cec4a0) * $signed(16'h0);
  assign T23057 = T23058 ? 2'h3 : 2'h0;
  assign T23058 = T23055[6'h2c:6'h2c];
  assign T23059 = $signed(T23060) / $signed(22'h100000);
  assign T23060 = $signed(31'h3f641b8d) * $signed(16'h1);
  assign T23061 = T18725[1'h0:1'h0];
  assign T23062 = T23077 ? twiddle4_1_47_real : twiddle4_1_46_real;
  assign twiddle4_1_46_real = T23068 + T23063;
  assign T23063 = {T23066, T23064};
  assign T23064 = $signed(T23065) / $signed(22'h100000);
  assign T23065 = $signed(29'h9008b6a) * $signed(16'h0);
  assign T23066 = T23067 ? 2'h3 : 2'h0;
  assign T23067 = T23064[6'h2c:6'h2c];
  assign T23068 = $signed(T23069) / $signed(22'h100000);
  assign T23069 = $signed(31'h3f5d1d1c) * $signed(16'h1);
  assign twiddle4_1_47_real = T23075 + T23070;
  assign T23070 = {T23073, T23071};
  assign T23071 = $signed(T23072) / $signed(22'h100000);
  assign T23072 = $signed(29'h9324ca6) * $signed(16'h0);
  assign T23073 = T23074 ? 2'h3 : 2'h0;
  assign T23074 = T23071[6'h2c:6'h2c];
  assign T23075 = $signed(T23076) / $signed(22'h100000);
  assign T23076 = $signed(31'h3f55f796) * $signed(16'h1);
  assign T23077 = T18725[1'h0:1'h0];
  assign T23078 = T18725[1'h1:1'h1];
  assign T23079 = T18725[2'h2:2'h2];
  assign T23080 = T18725[2'h3:2'h3];
  assign T23081 = T23222 ? T23152 : T23082;
  assign T23082 = T23151 ? T23117 : T23083;
  assign T23083 = T23116 ? T23100 : T23084;
  assign T23084 = T23099 ? twiddle4_1_49_real : twiddle4_1_48_real;
  assign twiddle4_1_48_real = T23090 + T23085;
  assign T23085 = {T23088, T23086};
  assign T23086 = $signed(T23087) / $signed(22'h100000);
  assign T23087 = $signed(29'h9640837) * $signed(16'h0);
  assign T23088 = T23089 ? 2'h3 : 2'h0;
  assign T23089 = T23086[6'h2c:6'h2c];
  assign T23090 = $signed(T23091) / $signed(22'h100000);
  assign T23091 = $signed(31'h3f4eaafe) * $signed(16'h1);
  assign twiddle4_1_49_real = T23097 + T23092;
  assign T23092 = {T23095, T23093};
  assign T23093 = $signed(T23094) / $signed(22'h100000);
  assign T23094 = $signed(29'h995bdfc) * $signed(16'h0);
  assign T23095 = T23096 ? 2'h3 : 2'h0;
  assign T23096 = T23093[6'h2c:6'h2c];
  assign T23097 = $signed(T23098) / $signed(22'h100000);
  assign T23098 = $signed(31'h3f473758) * $signed(16'h1);
  assign T23099 = T18725[1'h0:1'h0];
  assign T23100 = T23115 ? twiddle4_1_51_real : twiddle4_1_50_real;
  assign twiddle4_1_50_real = T23106 + T23101;
  assign T23101 = {T23104, T23102};
  assign T23102 = $signed(T23103) / $signed(22'h100000);
  assign T23103 = $signed(29'h9c76dd8) * $signed(16'h0);
  assign T23104 = T23105 ? 2'h3 : 2'h0;
  assign T23105 = T23102[6'h2c:6'h2c];
  assign T23106 = $signed(T23107) / $signed(22'h100000);
  assign T23107 = $signed(31'h3f3f9cab) * $signed(16'h1);
  assign twiddle4_1_51_real = T23113 + T23108;
  assign T23108 = {T23111, T23109};
  assign T23109 = $signed(T23110) / $signed(22'h100000);
  assign T23110 = $signed(29'h9f917ab) * $signed(16'h0);
  assign T23111 = T23112 ? 2'h3 : 2'h0;
  assign T23112 = T23109[6'h2c:6'h2c];
  assign T23113 = $signed(T23114) / $signed(22'h100000);
  assign T23114 = $signed(31'h3f37daf9) * $signed(16'h1);
  assign T23115 = T18725[1'h0:1'h0];
  assign T23116 = T18725[1'h1:1'h1];
  assign T23117 = T23150 ? T23134 : T23118;
  assign T23118 = T23133 ? twiddle4_1_53_real : twiddle4_1_52_real;
  assign twiddle4_1_52_real = T23124 + T23119;
  assign T23119 = {T23122, T23120};
  assign T23120 = $signed(T23121) / $signed(22'h100000);
  assign T23121 = $signed(29'ha2abb58) * $signed(16'h0);
  assign T23122 = T23123 ? 2'h3 : 2'h0;
  assign T23123 = T23120[6'h2c:6'h2c];
  assign T23124 = $signed(T23125) / $signed(22'h100000);
  assign T23125 = $signed(31'h3f2ff249) * $signed(16'h1);
  assign twiddle4_1_53_real = T23131 + T23126;
  assign T23126 = {T23129, T23127};
  assign T23127 = $signed(T23128) / $signed(22'h100000);
  assign T23128 = $signed(29'ha5c58bf) * $signed(16'h0);
  assign T23129 = T23130 ? 2'h3 : 2'h0;
  assign T23130 = T23127[6'h2c:6'h2c];
  assign T23131 = $signed(T23132) / $signed(22'h100000);
  assign T23132 = $signed(31'h3f27e29f) * $signed(16'h1);
  assign T23133 = T18725[1'h0:1'h0];
  assign T23134 = T23149 ? twiddle4_1_55_real : twiddle4_1_54_real;
  assign twiddle4_1_54_real = T23140 + T23135;
  assign T23135 = {T23138, T23136};
  assign T23136 = $signed(T23137) / $signed(22'h100000);
  assign T23137 = $signed(29'ha8defc2) * $signed(16'h0);
  assign T23138 = T23139 ? 2'h3 : 2'h0;
  assign T23139 = T23136[6'h2c:6'h2c];
  assign T23140 = $signed(T23141) / $signed(22'h100000);
  assign T23141 = $signed(31'h3f1fabff) * $signed(16'h1);
  assign twiddle4_1_55_real = T23147 + T23142;
  assign T23142 = {T23145, T23143};
  assign T23143 = $signed(T23144) / $signed(22'h100000);
  assign T23144 = $signed(29'habf8043) * $signed(16'h0);
  assign T23145 = T23146 ? 2'h3 : 2'h0;
  assign T23146 = T23143[6'h2c:6'h2c];
  assign T23147 = $signed(T23148) / $signed(22'h100000);
  assign T23148 = $signed(31'h3f174e6f) * $signed(16'h1);
  assign T23149 = T18725[1'h0:1'h0];
  assign T23150 = T18725[1'h1:1'h1];
  assign T23151 = T18725[2'h2:2'h2];
  assign T23152 = T23221 ? T23187 : T23153;
  assign T23153 = T23186 ? T23170 : T23154;
  assign T23154 = T23169 ? twiddle4_1_57_real : twiddle4_1_56_real;
  assign twiddle4_1_56_real = T23160 + T23155;
  assign T23155 = {T23158, T23156};
  assign T23156 = $signed(T23157) / $signed(22'h100000);
  assign T23157 = $signed(29'haf10a22) * $signed(16'h0);
  assign T23158 = T23159 ? 2'h3 : 2'h0;
  assign T23159 = T23156[6'h2c:6'h2c];
  assign T23160 = $signed(T23161) / $signed(22'h100000);
  assign T23161 = $signed(31'h3f0ec9f4) * $signed(16'h1);
  assign twiddle4_1_57_real = T23167 + T23162;
  assign T23162 = {T23165, T23163};
  assign T23163 = $signed(T23164) / $signed(22'h100000);
  assign T23164 = $signed(29'hb228d41) * $signed(16'h0);
  assign T23165 = T23166 ? 2'h3 : 2'h0;
  assign T23166 = T23163[6'h2c:6'h2c];
  assign T23167 = $signed(T23168) / $signed(22'h100000);
  assign T23168 = $signed(31'h3f061e94) * $signed(16'h1);
  assign T23169 = T18725[1'h0:1'h0];
  assign T23170 = T23185 ? twiddle4_1_59_real : twiddle4_1_58_real;
  assign twiddle4_1_58_real = T23176 + T23171;
  assign T23171 = {T23174, T23172};
  assign T23172 = $signed(T23173) / $signed(22'h100000);
  assign T23173 = $signed(29'hb540982) * $signed(16'h0);
  assign T23174 = T23175 ? 2'h3 : 2'h0;
  assign T23175 = T23172[6'h2c:6'h2c];
  assign T23176 = $signed(T23177) / $signed(22'h100000);
  assign T23177 = $signed(31'h3efd4c53) * $signed(16'h1);
  assign twiddle4_1_59_real = T23183 + T23178;
  assign T23178 = {T23181, T23179};
  assign T23179 = $signed(T23180) / $signed(22'h100000);
  assign T23180 = $signed(29'hb857ec6) * $signed(16'h0);
  assign T23181 = T23182 ? 2'h3 : 2'h0;
  assign T23182 = T23179[6'h2c:6'h2c];
  assign T23183 = $signed(T23184) / $signed(22'h100000);
  assign T23184 = $signed(31'h3ef45338) * $signed(16'h1);
  assign T23185 = T18725[1'h0:1'h0];
  assign T23186 = T18725[1'h1:1'h1];
  assign T23187 = T23220 ? T23204 : T23188;
  assign T23188 = T23203 ? twiddle4_1_61_real : twiddle4_1_60_real;
  assign twiddle4_1_60_real = T23194 + T23189;
  assign T23189 = {T23192, T23190};
  assign T23190 = $signed(T23191) / $signed(22'h100000);
  assign T23191 = $signed(29'hbb6ecef) * $signed(16'h0);
  assign T23192 = T23193 ? 2'h3 : 2'h0;
  assign T23193 = T23190[6'h2c:6'h2c];
  assign T23194 = $signed(T23195) / $signed(22'h100000);
  assign T23195 = $signed(31'h3eeb3347) * $signed(16'h1);
  assign twiddle4_1_61_real = T23201 + T23196;
  assign T23196 = {T23199, T23197};
  assign T23197 = $signed(T23198) / $signed(22'h100000);
  assign T23198 = $signed(29'hbe853dd) * $signed(16'h0);
  assign T23199 = T23200 ? 2'h3 : 2'h0;
  assign T23200 = T23197[6'h2c:6'h2c];
  assign T23201 = $signed(T23202) / $signed(22'h100000);
  assign T23202 = $signed(31'h3ee1ec86) * $signed(16'h1);
  assign T23203 = T18725[1'h0:1'h0];
  assign T23204 = T23219 ? twiddle4_1_63_real : twiddle4_1_62_real;
  assign twiddle4_1_62_real = T23210 + T23205;
  assign T23205 = {T23208, T23206};
  assign T23206 = $signed(T23207) / $signed(22'h100000);
  assign T23207 = $signed(29'hc19b374) * $signed(16'h0);
  assign T23208 = T23209 ? 2'h3 : 2'h0;
  assign T23209 = T23206[6'h2c:6'h2c];
  assign T23210 = $signed(T23211) / $signed(22'h100000);
  assign T23211 = $signed(31'h3ed87efb) * $signed(16'h1);
  assign twiddle4_1_63_real = T23217 + T23212;
  assign T23212 = {T23215, T23213};
  assign T23213 = $signed(T23214) / $signed(22'h100000);
  assign T23214 = $signed(29'hc4b0b93) * $signed(16'h0);
  assign T23215 = T23216 ? 2'h3 : 2'h0;
  assign T23216 = T23213[6'h2c:6'h2c];
  assign T23217 = $signed(T23218) / $signed(22'h100000);
  assign T23218 = $signed(31'h3eceeaad) * $signed(16'h1);
  assign T23219 = T18725[1'h0:1'h0];
  assign T23220 = T18725[1'h1:1'h1];
  assign T23221 = T18725[2'h2:2'h2];
  assign T23222 = T18725[2'h3:2'h3];
  assign T23223 = T18725[3'h4:3'h4];
  assign T23224 = T22938[6'h2e:6'h2e];
  assign T23225 = T18725[3'h5:3'h5];
  assign T23226 = {T23756, T23227};
  assign T23227 = T23755 ? T23501 : T23228;
  assign T23228 = T23500 ? T23371 : T23229;
  assign T23229 = T23370 ? T23300 : T23230;
  assign T23230 = T23299 ? T23265 : T23231;
  assign T23231 = T23264 ? T23248 : T23232;
  assign T23232 = T23247 ? twiddle4_1_65_real : twiddle4_1_64_real;
  assign twiddle4_1_64_real = T23238 + T23233;
  assign T23233 = {T23236, T23234};
  assign T23234 = $signed(T23235) / $signed(22'h100000);
  assign T23235 = $signed(29'hc7c5c1e) * $signed(16'h0);
  assign T23236 = T23237 ? 2'h3 : 2'h0;
  assign T23237 = T23234[6'h2c:6'h2c];
  assign T23238 = $signed(T23239) / $signed(22'h100000);
  assign T23239 = $signed(31'h3ec52f9f) * $signed(16'h1);
  assign twiddle4_1_65_real = T23245 + T23240;
  assign T23240 = {T23243, T23241};
  assign T23241 = $signed(T23242) / $signed(22'h100000);
  assign T23242 = $signed(29'hcada4f4) * $signed(16'h0);
  assign T23243 = T23244 ? 2'h3 : 2'h0;
  assign T23244 = T23241[6'h2c:6'h2c];
  assign T23245 = $signed(T23246) / $signed(22'h100000);
  assign T23246 = $signed(31'h3ebb4dda) * $signed(16'h1);
  assign T23247 = T18725[1'h0:1'h0];
  assign T23248 = T23263 ? twiddle4_1_67_real : twiddle4_1_66_real;
  assign twiddle4_1_66_real = T23254 + T23249;
  assign T23249 = {T23252, T23250};
  assign T23250 = $signed(T23251) / $signed(22'h100000);
  assign T23251 = $signed(29'hcdee5f9) * $signed(16'h0);
  assign T23252 = T23253 ? 2'h3 : 2'h0;
  assign T23253 = T23250[6'h2c:6'h2c];
  assign T23254 = $signed(T23255) / $signed(22'h100000);
  assign T23255 = $signed(31'h3eb14562) * $signed(16'h1);
  assign twiddle4_1_67_real = T23261 + T23256;
  assign T23256 = {T23259, T23257};
  assign T23257 = $signed(T23258) / $signed(22'h100000);
  assign T23258 = $signed(29'hd101f0d) * $signed(16'h0);
  assign T23259 = T23260 ? 2'h3 : 2'h0;
  assign T23260 = T23257[6'h2c:6'h2c];
  assign T23261 = $signed(T23262) / $signed(22'h100000);
  assign T23262 = $signed(31'h3ea7163f) * $signed(16'h1);
  assign T23263 = T18725[1'h0:1'h0];
  assign T23264 = T18725[1'h1:1'h1];
  assign T23265 = T23298 ? T23282 : T23266;
  assign T23266 = T23281 ? twiddle4_1_69_real : twiddle4_1_68_real;
  assign twiddle4_1_68_real = T23272 + T23267;
  assign T23267 = {T23270, T23268};
  assign T23268 = $signed(T23269) / $signed(22'h100000);
  assign T23269 = $signed(29'hd415012) * $signed(16'h0);
  assign T23270 = T23271 ? 2'h3 : 2'h0;
  assign T23271 = T23268[6'h2c:6'h2c];
  assign T23272 = $signed(T23273) / $signed(22'h100000);
  assign T23273 = $signed(31'h3e9cc076) * $signed(16'h1);
  assign twiddle4_1_69_real = T23279 + T23274;
  assign T23274 = {T23277, T23275};
  assign T23275 = $signed(T23276) / $signed(22'h100000);
  assign T23276 = $signed(29'hd7278ea) * $signed(16'h0);
  assign T23277 = T23278 ? 2'h3 : 2'h0;
  assign T23278 = T23275[6'h2c:6'h2c];
  assign T23279 = $signed(T23280) / $signed(22'h100000);
  assign T23280 = $signed(31'h3e92440d) * $signed(16'h1);
  assign T23281 = T18725[1'h0:1'h0];
  assign T23282 = T23297 ? twiddle4_1_71_real : twiddle4_1_70_real;
  assign twiddle4_1_70_real = T23288 + T23283;
  assign T23283 = {T23286, T23284};
  assign T23284 = $signed(T23285) / $signed(22'h100000);
  assign T23285 = $signed(29'hda39977) * $signed(16'h0);
  assign T23286 = T23287 ? 2'h3 : 2'h0;
  assign T23287 = T23284[6'h2c:6'h2c];
  assign T23288 = $signed(T23289) / $signed(22'h100000);
  assign T23289 = $signed(31'h3e87a10b) * $signed(16'h1);
  assign twiddle4_1_71_real = T23295 + T23290;
  assign T23290 = {T23293, T23291};
  assign T23291 = $signed(T23292) / $signed(22'h100000);
  assign T23292 = $signed(29'hdd4b19a) * $signed(16'h0);
  assign T23293 = T23294 ? 2'h3 : 2'h0;
  assign T23294 = T23291[6'h2c:6'h2c];
  assign T23295 = $signed(T23296) / $signed(22'h100000);
  assign T23296 = $signed(31'h3e7cd778) * $signed(16'h1);
  assign T23297 = T18725[1'h0:1'h0];
  assign T23298 = T18725[1'h1:1'h1];
  assign T23299 = T18725[2'h2:2'h2];
  assign T23300 = T23369 ? T23335 : T23301;
  assign T23301 = T23334 ? T23318 : T23302;
  assign T23302 = T23317 ? twiddle4_1_73_real : twiddle4_1_72_real;
  assign twiddle4_1_72_real = T23308 + T23303;
  assign T23303 = {T23306, T23304};
  assign T23304 = $signed(T23305) / $signed(22'h100000);
  assign T23305 = $signed(29'he05c135) * $signed(16'h0);
  assign T23306 = T23307 ? 2'h3 : 2'h0;
  assign T23307 = T23304[6'h2c:6'h2c];
  assign T23308 = $signed(T23309) / $signed(22'h100000);
  assign T23309 = $signed(31'h3e71e758) * $signed(16'h1);
  assign twiddle4_1_73_real = T23315 + T23310;
  assign T23310 = {T23313, T23311};
  assign T23311 = $signed(T23312) / $signed(22'h100000);
  assign T23312 = $signed(29'he36c829) * $signed(16'h0);
  assign T23313 = T23314 ? 2'h3 : 2'h0;
  assign T23314 = T23311[6'h2c:6'h2c];
  assign T23315 = $signed(T23316) / $signed(22'h100000);
  assign T23316 = $signed(31'h3e66d0b4) * $signed(16'h1);
  assign T23317 = T18725[1'h0:1'h0];
  assign T23318 = T23333 ? twiddle4_1_75_real : twiddle4_1_74_real;
  assign twiddle4_1_74_real = T23324 + T23319;
  assign T23319 = {T23322, T23320};
  assign T23320 = $signed(T23321) / $signed(22'h100000);
  assign T23321 = $signed(29'he67c659) * $signed(16'h0);
  assign T23322 = T23323 ? 2'h3 : 2'h0;
  assign T23323 = T23320[6'h2c:6'h2c];
  assign T23324 = $signed(T23325) / $signed(22'h100000);
  assign T23325 = $signed(31'h3e5b9392) * $signed(16'h1);
  assign twiddle4_1_75_real = T23331 + T23326;
  assign T23326 = {T23329, T23327};
  assign T23327 = $signed(T23328) / $signed(22'h100000);
  assign T23328 = $signed(29'he98bba6) * $signed(16'h0);
  assign T23329 = T23330 ? 2'h3 : 2'h0;
  assign T23330 = T23327[6'h2c:6'h2c];
  assign T23331 = $signed(T23332) / $signed(22'h100000);
  assign T23332 = $signed(31'h3e502ff8) * $signed(16'h1);
  assign T23333 = T18725[1'h0:1'h0];
  assign T23334 = T18725[1'h1:1'h1];
  assign T23335 = T23368 ? T23352 : T23336;
  assign T23336 = T23351 ? twiddle4_1_77_real : twiddle4_1_76_real;
  assign twiddle4_1_76_real = T23342 + T23337;
  assign T23337 = {T23340, T23338};
  assign T23338 = $signed(T23339) / $signed(22'h100000);
  assign T23339 = $signed(29'hec9a7f2) * $signed(16'h0);
  assign T23340 = T23341 ? 2'h3 : 2'h0;
  assign T23341 = T23338[6'h2c:6'h2c];
  assign T23342 = $signed(T23343) / $signed(22'h100000);
  assign T23343 = $signed(31'h3e44a5ee) * $signed(16'h1);
  assign twiddle4_1_77_real = T23349 + T23344;
  assign T23344 = {T23347, T23345};
  assign T23345 = $signed(T23346) / $signed(22'h100000);
  assign T23346 = $signed(29'hefa8b1f) * $signed(16'h0);
  assign T23347 = T23348 ? 2'h3 : 2'h0;
  assign T23348 = T23345[6'h2c:6'h2c];
  assign T23349 = $signed(T23350) / $signed(22'h100000);
  assign T23350 = $signed(31'h3e38f57c) * $signed(16'h1);
  assign T23351 = T18725[1'h0:1'h0];
  assign T23352 = T23367 ? twiddle4_1_79_real : twiddle4_1_78_real;
  assign twiddle4_1_78_real = T23358 + T23353;
  assign T23353 = {T23356, T23354};
  assign T23354 = $signed(T23355) / $signed(22'h100000);
  assign T23355 = $signed(29'hf2b650f) * $signed(16'h0);
  assign T23356 = T23357 ? 2'h3 : 2'h0;
  assign T23357 = T23354[6'h2c:6'h2c];
  assign T23358 = $signed(T23359) / $signed(22'h100000);
  assign T23359 = $signed(31'h3e2d1ea7) * $signed(16'h1);
  assign twiddle4_1_79_real = T23365 + T23360;
  assign T23360 = {T23363, T23361};
  assign T23361 = $signed(T23362) / $signed(22'h100000);
  assign T23362 = $signed(29'hf5c35a3) * $signed(16'h0);
  assign T23363 = T23364 ? 2'h3 : 2'h0;
  assign T23364 = T23361[6'h2c:6'h2c];
  assign T23365 = $signed(T23366) / $signed(22'h100000);
  assign T23366 = $signed(31'h3e212179) * $signed(16'h1);
  assign T23367 = T18725[1'h0:1'h0];
  assign T23368 = T18725[1'h1:1'h1];
  assign T23369 = T18725[2'h2:2'h2];
  assign T23370 = T18725[2'h3:2'h3];
  assign T23371 = T23499 ? T23437 : T23372;
  assign T23372 = T23436 ? T23406 : T23373;
  assign T23373 = T23405 ? T23390 : T23374;
  assign T23374 = T23389 ? twiddle4_1_81_real : twiddle4_1_80_real;
  assign twiddle4_1_80_real = T23380 + T23375;
  assign T23375 = {T23378, T23376};
  assign T23376 = $signed(T23377) / $signed(22'h100000);
  assign T23377 = $signed(29'hf8cfcbd) * $signed(16'h0);
  assign T23378 = T23379 ? 2'h3 : 2'h0;
  assign T23379 = T23376[6'h2c:6'h2c];
  assign T23380 = $signed(T23381) / $signed(22'h100000);
  assign T23381 = $signed(31'h3e14fdf7) * $signed(16'h1);
  assign twiddle4_1_81_real = T23387 + T23382;
  assign T23382 = {T23385, T23383};
  assign T23383 = $signed(T23384) / $signed(22'h100000);
  assign T23384 = $signed(29'hfbdba40) * $signed(16'h0);
  assign T23385 = T23386 ? 2'h3 : 2'h0;
  assign T23386 = T23383[6'h2c:6'h2c];
  assign T23387 = $signed(T23388) / $signed(22'h100000);
  assign T23388 = $signed(31'h3e08b429) * $signed(16'h1);
  assign T23389 = T18725[1'h0:1'h0];
  assign T23390 = T23404 ? twiddle4_1_83_real : twiddle4_1_82_real;
  assign twiddle4_1_82_real = T23396 + T23391;
  assign T23391 = {T23394, T23392};
  assign T23392 = $signed(T23393) / $signed(22'h100000);
  assign T23393 = $signed(29'hfee6e0d) * $signed(16'h0);
  assign T23394 = T23395 ? 2'h3 : 2'h0;
  assign T23395 = T23392[6'h2c:6'h2c];
  assign T23396 = $signed(T23397) / $signed(22'h100000);
  assign T23397 = $signed(31'h3dfc4418) * $signed(16'h1);
  assign twiddle4_1_83_real = T23402 + T23398;
  assign T23398 = {T23401, T23399};
  assign T23399 = $signed(T23400) / $signed(22'h100000);
  assign T23400 = $signed(30'h101f1806) * $signed(16'h0);
  assign T23401 = T23399[6'h2d:6'h2d];
  assign T23402 = $signed(T23403) / $signed(22'h100000);
  assign T23403 = $signed(31'h3defadca) * $signed(16'h1);
  assign T23404 = T18725[1'h0:1'h0];
  assign T23405 = T18725[1'h1:1'h1];
  assign T23406 = T23435 ? T23421 : T23407;
  assign T23407 = T23420 ? twiddle4_1_85_real : twiddle4_1_84_real;
  assign twiddle4_1_84_real = T23412 + T23408;
  assign T23408 = {T23411, T23409};
  assign T23409 = $signed(T23410) / $signed(22'h100000);
  assign T23410 = $signed(30'h104fb80e) * $signed(16'h0);
  assign T23411 = T23409[6'h2d:6'h2d];
  assign T23412 = $signed(T23413) / $signed(22'h100000);
  assign T23413 = $signed(31'h3de2f147) * $signed(16'h1);
  assign twiddle4_1_85_real = T23418 + T23414;
  assign T23414 = {T23417, T23415};
  assign T23415 = $signed(T23416) / $signed(22'h100000);
  assign T23416 = $signed(30'h10804e05) * $signed(16'h0);
  assign T23417 = T23415[6'h2d:6'h2d];
  assign T23418 = $signed(T23419) / $signed(22'h100000);
  assign T23419 = $signed(31'h3dd60e98) * $signed(16'h1);
  assign T23420 = T18725[1'h0:1'h0];
  assign T23421 = T23434 ? twiddle4_1_87_real : twiddle4_1_86_real;
  assign twiddle4_1_86_real = T23426 + T23422;
  assign T23422 = {T23425, T23423};
  assign T23423 = $signed(T23424) / $signed(22'h100000);
  assign T23424 = $signed(30'h10b0d9cf) * $signed(16'h0);
  assign T23425 = T23423[6'h2d:6'h2d];
  assign T23426 = $signed(T23427) / $signed(22'h100000);
  assign T23427 = $signed(31'h3dc905c4) * $signed(16'h1);
  assign twiddle4_1_87_real = T23432 + T23428;
  assign T23428 = {T23431, T23429};
  assign T23429 = $signed(T23430) / $signed(22'h100000);
  assign T23430 = $signed(30'h10e15b4e) * $signed(16'h0);
  assign T23431 = T23429[6'h2d:6'h2d];
  assign T23432 = $signed(T23433) / $signed(22'h100000);
  assign T23433 = $signed(31'h3dbbd6d4) * $signed(16'h1);
  assign T23434 = T18725[1'h0:1'h0];
  assign T23435 = T18725[1'h1:1'h1];
  assign T23436 = T18725[2'h2:2'h2];
  assign T23437 = T23498 ? T23468 : T23438;
  assign T23438 = T23467 ? T23453 : T23439;
  assign T23439 = T23452 ? twiddle4_1_89_real : twiddle4_1_88_real;
  assign twiddle4_1_88_real = T23444 + T23440;
  assign T23440 = {T23443, T23441};
  assign T23441 = $signed(T23442) / $signed(22'h100000);
  assign T23442 = $signed(30'h1111d262) * $signed(16'h0);
  assign T23443 = T23441[6'h2d:6'h2d];
  assign T23444 = $signed(T23445) / $signed(22'h100000);
  assign T23445 = $signed(31'h3dae81ce) * $signed(16'h1);
  assign twiddle4_1_89_real = T23450 + T23446;
  assign T23446 = {T23449, T23447};
  assign T23447 = $signed(T23448) / $signed(22'h100000);
  assign T23448 = $signed(30'h11423eef) * $signed(16'h0);
  assign T23449 = T23447[6'h2d:6'h2d];
  assign T23450 = $signed(T23451) / $signed(22'h100000);
  assign T23451 = $signed(31'h3da106bd) * $signed(16'h1);
  assign T23452 = T18725[1'h0:1'h0];
  assign T23453 = T23466 ? twiddle4_1_91_real : twiddle4_1_90_real;
  assign twiddle4_1_90_real = T23458 + T23454;
  assign T23454 = {T23457, T23455};
  assign T23455 = $signed(T23456) / $signed(22'h100000);
  assign T23456 = $signed(30'h1172a0d7) * $signed(16'h0);
  assign T23457 = T23455[6'h2d:6'h2d];
  assign T23458 = $signed(T23459) / $signed(22'h100000);
  assign T23459 = $signed(31'h3d9365a7) * $signed(16'h1);
  assign twiddle4_1_91_real = T23464 + T23460;
  assign T23460 = {T23463, T23461};
  assign T23461 = $signed(T23462) / $signed(22'h100000);
  assign T23462 = $signed(30'h11a2f7fb) * $signed(16'h0);
  assign T23463 = T23461[6'h2d:6'h2d];
  assign T23464 = $signed(T23465) / $signed(22'h100000);
  assign T23465 = $signed(31'h3d859e96) * $signed(16'h1);
  assign T23466 = T18725[1'h0:1'h0];
  assign T23467 = T18725[1'h1:1'h1];
  assign T23468 = T23497 ? T23483 : T23469;
  assign T23469 = T23482 ? twiddle4_1_93_real : twiddle4_1_92_real;
  assign twiddle4_1_92_real = T23474 + T23470;
  assign T23470 = {T23473, T23471};
  assign T23471 = $signed(T23472) / $signed(22'h100000);
  assign T23472 = $signed(30'h11d3443f) * $signed(16'h0);
  assign T23473 = T23471[6'h2d:6'h2d];
  assign T23474 = $signed(T23475) / $signed(22'h100000);
  assign T23475 = $signed(31'h3d77b191) * $signed(16'h1);
  assign twiddle4_1_93_real = T23480 + T23476;
  assign T23476 = {T23479, T23477};
  assign T23477 = $signed(T23478) / $signed(22'h100000);
  assign T23478 = $signed(30'h12038583) * $signed(16'h0);
  assign T23479 = T23477[6'h2d:6'h2d];
  assign T23480 = $signed(T23481) / $signed(22'h100000);
  assign T23481 = $signed(31'h3d699ea2) * $signed(16'h1);
  assign T23482 = T18725[1'h0:1'h0];
  assign T23483 = T23496 ? twiddle4_1_95_real : twiddle4_1_94_real;
  assign twiddle4_1_94_real = T23488 + T23484;
  assign T23484 = {T23487, T23485};
  assign T23485 = $signed(T23486) / $signed(22'h100000);
  assign T23486 = $signed(30'h1233bbab) * $signed(16'h0);
  assign T23487 = T23485[6'h2d:6'h2d];
  assign T23488 = $signed(T23489) / $signed(22'h100000);
  assign T23489 = $signed(31'h3d5b65d1) * $signed(16'h1);
  assign twiddle4_1_95_real = T23494 + T23490;
  assign T23490 = {T23493, T23491};
  assign T23491 = $signed(T23492) / $signed(22'h100000);
  assign T23492 = $signed(30'h1263e699) * $signed(16'h0);
  assign T23493 = T23491[6'h2d:6'h2d];
  assign T23494 = $signed(T23495) / $signed(22'h100000);
  assign T23495 = $signed(31'h3d4d0727) * $signed(16'h1);
  assign T23496 = T18725[1'h0:1'h0];
  assign T23497 = T18725[1'h1:1'h1];
  assign T23498 = T18725[2'h2:2'h2];
  assign T23499 = T18725[2'h3:2'h3];
  assign T23500 = T18725[3'h4:3'h4];
  assign T23501 = T23754 ? T23628 : T23502;
  assign T23502 = T23627 ? T23565 : T23503;
  assign T23503 = T23564 ? T23534 : T23504;
  assign T23504 = T23533 ? T23519 : T23505;
  assign T23505 = T23518 ? twiddle4_1_97_real : twiddle4_1_96_real;
  assign twiddle4_1_96_real = T23510 + T23506;
  assign T23506 = {T23509, T23507};
  assign T23507 = $signed(T23508) / $signed(22'h100000);
  assign T23508 = $signed(30'h1294062e) * $signed(16'h0);
  assign T23509 = T23507[6'h2d:6'h2d];
  assign T23510 = $signed(T23511) / $signed(22'h100000);
  assign T23511 = $signed(31'h3d3e82ad) * $signed(16'h1);
  assign twiddle4_1_97_real = T23516 + T23512;
  assign T23512 = {T23515, T23513};
  assign T23513 = $signed(T23514) / $signed(22'h100000);
  assign T23514 = $signed(30'h12c41a4e) * $signed(16'h0);
  assign T23515 = T23513[6'h2d:6'h2d];
  assign T23516 = $signed(T23517) / $signed(22'h100000);
  assign T23517 = $signed(31'h3d2fd86c) * $signed(16'h1);
  assign T23518 = T18725[1'h0:1'h0];
  assign T23519 = T23532 ? twiddle4_1_99_real : twiddle4_1_98_real;
  assign twiddle4_1_98_real = T23524 + T23520;
  assign T23520 = {T23523, T23521};
  assign T23521 = $signed(T23522) / $signed(22'h100000);
  assign T23522 = $signed(30'h12f422da) * $signed(16'h0);
  assign T23523 = T23521[6'h2d:6'h2d];
  assign T23524 = $signed(T23525) / $signed(22'h100000);
  assign T23525 = $signed(31'h3d21086c) * $signed(16'h1);
  assign twiddle4_1_99_real = T23530 + T23526;
  assign T23526 = {T23529, T23527};
  assign T23527 = $signed(T23528) / $signed(22'h100000);
  assign T23528 = $signed(30'h13241fb6) * $signed(16'h0);
  assign T23529 = T23527[6'h2d:6'h2d];
  assign T23530 = $signed(T23531) / $signed(22'h100000);
  assign T23531 = $signed(31'h3d1212b7) * $signed(16'h1);
  assign T23532 = T18725[1'h0:1'h0];
  assign T23533 = T18725[1'h1:1'h1];
  assign T23534 = T23563 ? T23549 : T23535;
  assign T23535 = T23548 ? twiddle4_1_101_real : twiddle4_1_100_real;
  assign twiddle4_1_100_real = T23540 + T23536;
  assign T23536 = {T23539, T23537};
  assign T23537 = $signed(T23538) / $signed(22'h100000);
  assign T23538 = $signed(30'h135410c2) * $signed(16'h0);
  assign T23539 = T23537[6'h2d:6'h2d];
  assign T23540 = $signed(T23541) / $signed(22'h100000);
  assign T23541 = $signed(31'h3d02f756) * $signed(16'h1);
  assign twiddle4_1_101_real = T23546 + T23542;
  assign T23542 = {T23545, T23543};
  assign T23543 = $signed(T23544) / $signed(22'h100000);
  assign T23544 = $signed(30'h1383f5e3) * $signed(16'h0);
  assign T23545 = T23543[6'h2d:6'h2d];
  assign T23546 = $signed(T23547) / $signed(22'h100000);
  assign T23547 = $signed(31'h3cf3b653) * $signed(16'h1);
  assign T23548 = T18725[1'h0:1'h0];
  assign T23549 = T23562 ? twiddle4_1_103_real : twiddle4_1_102_real;
  assign twiddle4_1_102_real = T23554 + T23550;
  assign T23550 = {T23553, T23551};
  assign T23551 = $signed(T23552) / $signed(22'h100000);
  assign T23552 = $signed(30'h13b3cefa) * $signed(16'h0);
  assign T23553 = T23551[6'h2d:6'h2d];
  assign T23554 = $signed(T23555) / $signed(22'h100000);
  assign T23555 = $signed(31'h3ce44fb6) * $signed(16'h1);
  assign twiddle4_1_103_real = T23560 + T23556;
  assign T23556 = {T23559, T23557};
  assign T23557 = $signed(T23558) / $signed(22'h100000);
  assign T23558 = $signed(30'h13e39be9) * $signed(16'h0);
  assign T23559 = T23557[6'h2d:6'h2d];
  assign T23560 = $signed(T23561) / $signed(22'h100000);
  assign T23561 = $signed(31'h3cd4c38a) * $signed(16'h1);
  assign T23562 = T18725[1'h0:1'h0];
  assign T23563 = T18725[1'h1:1'h1];
  assign T23564 = T18725[2'h2:2'h2];
  assign T23565 = T23626 ? T23596 : T23566;
  assign T23566 = T23595 ? T23581 : T23567;
  assign T23567 = T23580 ? twiddle4_1_105_real : twiddle4_1_104_real;
  assign twiddle4_1_104_real = T23572 + T23568;
  assign T23568 = {T23571, T23569};
  assign T23569 = $signed(T23570) / $signed(22'h100000);
  assign T23570 = $signed(30'h14135c94) * $signed(16'h0);
  assign T23571 = T23569[6'h2d:6'h2d];
  assign T23572 = $signed(T23573) / $signed(22'h100000);
  assign T23573 = $signed(31'h3cc511d8) * $signed(16'h1);
  assign twiddle4_1_105_real = T23578 + T23574;
  assign T23574 = {T23577, T23575};
  assign T23575 = $signed(T23576) / $signed(22'h100000);
  assign T23576 = $signed(30'h144310dc) * $signed(16'h0);
  assign T23577 = T23575[6'h2d:6'h2d];
  assign T23578 = $signed(T23579) / $signed(22'h100000);
  assign T23579 = $signed(31'h3cb53aaa) * $signed(16'h1);
  assign T23580 = T18725[1'h0:1'h0];
  assign T23581 = T23594 ? twiddle4_1_107_real : twiddle4_1_106_real;
  assign twiddle4_1_106_real = T23586 + T23582;
  assign T23582 = {T23585, T23583};
  assign T23583 = $signed(T23584) / $signed(22'h100000);
  assign T23584 = $signed(30'h1472b8a5) * $signed(16'h0);
  assign T23585 = T23583[6'h2d:6'h2d];
  assign T23586 = $signed(T23587) / $signed(22'h100000);
  assign T23587 = $signed(31'h3ca53e08) * $signed(16'h1);
  assign twiddle4_1_107_real = T23592 + T23588;
  assign T23588 = {T23591, T23589};
  assign T23589 = $signed(T23590) / $signed(22'h100000);
  assign T23590 = $signed(30'h14a253d1) * $signed(16'h0);
  assign T23591 = T23589[6'h2d:6'h2d];
  assign T23592 = $signed(T23593) / $signed(22'h100000);
  assign T23593 = $signed(31'h3c951bff) * $signed(16'h1);
  assign T23594 = T18725[1'h0:1'h0];
  assign T23595 = T18725[1'h1:1'h1];
  assign T23596 = T23625 ? T23611 : T23597;
  assign T23597 = T23610 ? twiddle4_1_109_real : twiddle4_1_108_real;
  assign twiddle4_1_108_real = T23602 + T23598;
  assign T23598 = {T23601, T23599};
  assign T23599 = $signed(T23600) / $signed(22'h100000);
  assign T23600 = $signed(30'h14d1e242) * $signed(16'h0);
  assign T23601 = T23599[6'h2d:6'h2d];
  assign T23602 = $signed(T23603) / $signed(22'h100000);
  assign T23603 = $signed(31'h3c84d496) * $signed(16'h1);
  assign twiddle4_1_109_real = T23608 + T23604;
  assign T23604 = {T23607, T23605};
  assign T23605 = $signed(T23606) / $signed(22'h100000);
  assign T23606 = $signed(30'h150163dc) * $signed(16'h0);
  assign T23607 = T23605[6'h2d:6'h2d];
  assign T23608 = $signed(T23609) / $signed(22'h100000);
  assign T23609 = $signed(31'h3c7467d8) * $signed(16'h1);
  assign T23610 = T18725[1'h0:1'h0];
  assign T23611 = T23624 ? twiddle4_1_111_real : twiddle4_1_110_real;
  assign twiddle4_1_110_real = T23616 + T23612;
  assign T23612 = {T23615, T23613};
  assign T23613 = $signed(T23614) / $signed(22'h100000);
  assign T23614 = $signed(30'h1530d880) * $signed(16'h0);
  assign T23615 = T23613[6'h2d:6'h2d];
  assign T23616 = $signed(T23617) / $signed(22'h100000);
  assign T23617 = $signed(31'h3c63d5d0) * $signed(16'h1);
  assign twiddle4_1_111_real = T23622 + T23618;
  assign T23618 = {T23621, T23619};
  assign T23619 = $signed(T23620) / $signed(22'h100000);
  assign T23620 = $signed(30'h15604012) * $signed(16'h0);
  assign T23621 = T23619[6'h2d:6'h2d];
  assign T23622 = $signed(T23623) / $signed(22'h100000);
  assign T23623 = $signed(31'h3c531e88) * $signed(16'h1);
  assign T23624 = T18725[1'h0:1'h0];
  assign T23625 = T18725[1'h1:1'h1];
  assign T23626 = T18725[2'h2:2'h2];
  assign T23627 = T18725[2'h3:2'h3];
  assign T23628 = T23753 ? T23691 : T23629;
  assign T23629 = T23690 ? T23660 : T23630;
  assign T23630 = T23659 ? T23645 : T23631;
  assign T23631 = T23644 ? twiddle4_1_113_real : twiddle4_1_112_real;
  assign twiddle4_1_112_real = T23636 + T23632;
  assign T23632 = {T23635, T23633};
  assign T23633 = $signed(T23634) / $signed(22'h100000);
  assign T23634 = $signed(30'h158f9a75) * $signed(16'h0);
  assign T23635 = T23633[6'h2d:6'h2d];
  assign T23636 = $signed(T23637) / $signed(22'h100000);
  assign T23637 = $signed(31'h3c424209) * $signed(16'h1);
  assign twiddle4_1_113_real = T23642 + T23638;
  assign T23638 = {T23641, T23639};
  assign T23639 = $signed(T23640) / $signed(22'h100000);
  assign T23640 = $signed(30'h15bee78b) * $signed(16'h0);
  assign T23641 = T23639[6'h2d:6'h2d];
  assign T23642 = $signed(T23643) / $signed(22'h100000);
  assign T23643 = $signed(31'h3c31405f) * $signed(16'h1);
  assign T23644 = T18725[1'h0:1'h0];
  assign T23645 = T23658 ? twiddle4_1_115_real : twiddle4_1_114_real;
  assign twiddle4_1_114_real = T23650 + T23646;
  assign T23646 = {T23649, T23647};
  assign T23647 = $signed(T23648) / $signed(22'h100000);
  assign T23648 = $signed(30'h15ee2737) * $signed(16'h0);
  assign T23649 = T23647[6'h2d:6'h2d];
  assign T23650 = $signed(T23651) / $signed(22'h100000);
  assign T23651 = $signed(31'h3c201994) * $signed(16'h1);
  assign twiddle4_1_115_real = T23656 + T23652;
  assign T23652 = {T23655, T23653};
  assign T23653 = $signed(T23654) / $signed(22'h100000);
  assign T23654 = $signed(30'h161d595c) * $signed(16'h0);
  assign T23655 = T23653[6'h2d:6'h2d];
  assign T23656 = $signed(T23657) / $signed(22'h100000);
  assign T23657 = $signed(31'h3c0ecdb2) * $signed(16'h1);
  assign T23658 = T18725[1'h0:1'h0];
  assign T23659 = T18725[1'h1:1'h1];
  assign T23660 = T23689 ? T23675 : T23661;
  assign T23661 = T23674 ? twiddle4_1_117_real : twiddle4_1_116_real;
  assign twiddle4_1_116_real = T23666 + T23662;
  assign T23662 = {T23665, T23663};
  assign T23663 = $signed(T23664) / $signed(22'h100000);
  assign T23664 = $signed(30'h164c7ddd) * $signed(16'h0);
  assign T23665 = T23663[6'h2d:6'h2d];
  assign T23666 = $signed(T23667) / $signed(22'h100000);
  assign T23667 = $signed(31'h3bfd5cc4) * $signed(16'h1);
  assign twiddle4_1_117_real = T23672 + T23668;
  assign T23668 = {T23671, T23669};
  assign T23669 = $signed(T23670) / $signed(22'h100000);
  assign T23670 = $signed(30'h167b949c) * $signed(16'h0);
  assign T23671 = T23669[6'h2d:6'h2d];
  assign T23672 = $signed(T23673) / $signed(22'h100000);
  assign T23673 = $signed(31'h3bebc6d5) * $signed(16'h1);
  assign T23674 = T18725[1'h0:1'h0];
  assign T23675 = T23688 ? twiddle4_1_119_real : twiddle4_1_118_real;
  assign twiddle4_1_118_real = T23680 + T23676;
  assign T23676 = {T23679, T23677};
  assign T23677 = $signed(T23678) / $signed(22'h100000);
  assign T23678 = $signed(30'h16aa9d7d) * $signed(16'h0);
  assign T23679 = T23677[6'h2d:6'h2d];
  assign T23680 = $signed(T23681) / $signed(22'h100000);
  assign T23681 = $signed(31'h3bda0bef) * $signed(16'h1);
  assign twiddle4_1_119_real = T23686 + T23682;
  assign T23682 = {T23685, T23683};
  assign T23683 = $signed(T23684) / $signed(22'h100000);
  assign T23684 = $signed(30'h16d99863) * $signed(16'h0);
  assign T23685 = T23683[6'h2d:6'h2d];
  assign T23686 = $signed(T23687) / $signed(22'h100000);
  assign T23687 = $signed(31'h3bc82c1e) * $signed(16'h1);
  assign T23688 = T18725[1'h0:1'h0];
  assign T23689 = T18725[1'h1:1'h1];
  assign T23690 = T18725[2'h2:2'h2];
  assign T23691 = T23752 ? T23722 : T23692;
  assign T23692 = T23721 ? T23707 : T23693;
  assign T23693 = T23706 ? twiddle4_1_121_real : twiddle4_1_120_real;
  assign twiddle4_1_120_real = T23698 + T23694;
  assign T23694 = {T23697, T23695};
  assign T23695 = $signed(T23696) / $signed(22'h100000);
  assign T23696 = $signed(30'h17088530) * $signed(16'h0);
  assign T23697 = T23695[6'h2d:6'h2d];
  assign T23698 = $signed(T23699) / $signed(22'h100000);
  assign T23699 = $signed(31'h3bb6276d) * $signed(16'h1);
  assign twiddle4_1_121_real = T23704 + T23700;
  assign T23700 = {T23703, T23701};
  assign T23701 = $signed(T23702) / $signed(22'h100000);
  assign T23702 = $signed(30'h173763c9) * $signed(16'h0);
  assign T23703 = T23701[6'h2d:6'h2d];
  assign T23704 = $signed(T23705) / $signed(22'h100000);
  assign T23705 = $signed(31'h3ba3fde7) * $signed(16'h1);
  assign T23706 = T18725[1'h0:1'h0];
  assign T23707 = T23720 ? twiddle4_1_123_real : twiddle4_1_122_real;
  assign twiddle4_1_122_real = T23712 + T23708;
  assign T23708 = {T23711, T23709};
  assign T23709 = $signed(T23710) / $signed(22'h100000);
  assign T23710 = $signed(30'h1766340f) * $signed(16'h0);
  assign T23711 = T23709[6'h2d:6'h2d];
  assign T23712 = $signed(T23713) / $signed(22'h100000);
  assign T23713 = $signed(31'h3b91af96) * $signed(16'h1);
  assign twiddle4_1_123_real = T23718 + T23714;
  assign T23714 = {T23717, T23715};
  assign T23715 = $signed(T23716) / $signed(22'h100000);
  assign T23716 = $signed(30'h1794f5e6) * $signed(16'h0);
  assign T23717 = T23715[6'h2d:6'h2d];
  assign T23718 = $signed(T23719) / $signed(22'h100000);
  assign T23719 = $signed(31'h3b7f3c87) * $signed(16'h1);
  assign T23720 = T18725[1'h0:1'h0];
  assign T23721 = T18725[1'h1:1'h1];
  assign T23722 = T23751 ? T23737 : T23723;
  assign T23723 = T23736 ? twiddle4_1_125_real : twiddle4_1_124_real;
  assign twiddle4_1_124_real = T23728 + T23724;
  assign T23724 = {T23727, T23725};
  assign T23725 = $signed(T23726) / $signed(22'h100000);
  assign T23726 = $signed(30'h17c3a931) * $signed(16'h0);
  assign T23727 = T23725[6'h2d:6'h2d];
  assign T23728 = $signed(T23729) / $signed(22'h100000);
  assign T23729 = $signed(31'h3b6ca4c4) * $signed(16'h1);
  assign twiddle4_1_125_real = T23734 + T23730;
  assign T23730 = {T23733, T23731};
  assign T23731 = $signed(T23732) / $signed(22'h100000);
  assign T23732 = $signed(30'h17f24dd3) * $signed(16'h0);
  assign T23733 = T23731[6'h2d:6'h2d];
  assign T23734 = $signed(T23735) / $signed(22'h100000);
  assign T23735 = $signed(31'h3b59e859) * $signed(16'h1);
  assign T23736 = T18725[1'h0:1'h0];
  assign T23737 = T23750 ? twiddle4_1_127_real : twiddle4_1_126_real;
  assign twiddle4_1_126_real = T23742 + T23738;
  assign T23738 = {T23741, T23739};
  assign T23739 = $signed(T23740) / $signed(22'h100000);
  assign T23740 = $signed(30'h1820e3b0) * $signed(16'h0);
  assign T23741 = T23739[6'h2d:6'h2d];
  assign T23742 = $signed(T23743) / $signed(22'h100000);
  assign T23743 = $signed(31'h3b470752) * $signed(16'h1);
  assign twiddle4_1_127_real = T23748 + T23744;
  assign T23744 = {T23747, T23745};
  assign T23745 = $signed(T23746) / $signed(22'h100000);
  assign T23746 = $signed(30'h184f6aaa) * $signed(16'h0);
  assign T23747 = T23745[6'h2d:6'h2d];
  assign T23748 = $signed(T23749) / $signed(22'h100000);
  assign T23749 = $signed(31'h3b3401bb) * $signed(16'h1);
  assign T23750 = T18725[1'h0:1'h0];
  assign T23751 = T18725[1'h1:1'h1];
  assign T23752 = T18725[2'h2:2'h2];
  assign T23753 = T18725[2'h3:2'h3];
  assign T23754 = T18725[3'h4:3'h4];
  assign T23755 = T18725[3'h5:3'h5];
  assign T23756 = T23227[6'h2e:6'h2e];
  assign T23757 = T18725[3'h6:3'h6];
  assign T23758 = {T24611, T23759};
  assign T23759 = T24610 ? T24228 : T23760;
  assign T23760 = T24227 ? T24015 : T23761;
  assign T23761 = T24014 ? T23888 : T23762;
  assign T23762 = T23887 ? T23825 : T23763;
  assign T23763 = T23824 ? T23794 : T23764;
  assign T23764 = T23793 ? T23779 : T23765;
  assign T23765 = T23778 ? twiddle4_1_129_real : twiddle4_1_128_real;
  assign twiddle4_1_128_real = T23770 + T23766;
  assign T23766 = {T23769, T23767};
  assign T23767 = $signed(T23768) / $signed(22'h100000);
  assign T23768 = $signed(30'h187de2a6) * $signed(16'h0);
  assign T23769 = T23767[6'h2d:6'h2d];
  assign T23770 = $signed(T23771) / $signed(22'h100000);
  assign T23771 = $signed(31'h3b20d79e) * $signed(16'h1);
  assign twiddle4_1_129_real = T23776 + T23772;
  assign T23772 = {T23775, T23773};
  assign T23773 = $signed(T23774) / $signed(22'h100000);
  assign T23774 = $signed(30'h18ac4b86) * $signed(16'h0);
  assign T23775 = T23773[6'h2d:6'h2d];
  assign T23776 = $signed(T23777) / $signed(22'h100000);
  assign T23777 = $signed(31'h3b0d8908) * $signed(16'h1);
  assign T23778 = T18725[1'h0:1'h0];
  assign T23779 = T23792 ? twiddle4_1_131_real : twiddle4_1_130_real;
  assign twiddle4_1_130_real = T23784 + T23780;
  assign T23780 = {T23783, T23781};
  assign T23781 = $signed(T23782) / $signed(22'h100000);
  assign T23782 = $signed(30'h18daa52e) * $signed(16'h0);
  assign T23783 = T23781[6'h2d:6'h2d];
  assign T23784 = $signed(T23785) / $signed(22'h100000);
  assign T23785 = $signed(31'h3afa1605) * $signed(16'h1);
  assign twiddle4_1_131_real = T23790 + T23786;
  assign T23786 = {T23789, T23787};
  assign T23787 = $signed(T23788) / $signed(22'h100000);
  assign T23788 = $signed(30'h1908ef81) * $signed(16'h0);
  assign T23789 = T23787[6'h2d:6'h2d];
  assign T23790 = $signed(T23791) / $signed(22'h100000);
  assign T23791 = $signed(31'h3ae67ea1) * $signed(16'h1);
  assign T23792 = T18725[1'h0:1'h0];
  assign T23793 = T18725[1'h1:1'h1];
  assign T23794 = T23823 ? T23809 : T23795;
  assign T23795 = T23808 ? twiddle4_1_133_real : twiddle4_1_132_real;
  assign twiddle4_1_132_real = T23800 + T23796;
  assign T23796 = {T23799, T23797};
  assign T23797 = $signed(T23798) / $signed(22'h100000);
  assign T23798 = $signed(30'h19372a63) * $signed(16'h0);
  assign T23799 = T23797[6'h2d:6'h2d];
  assign T23800 = $signed(T23801) / $signed(22'h100000);
  assign T23801 = $signed(31'h3ad2c2e7) * $signed(16'h1);
  assign twiddle4_1_133_real = T23806 + T23802;
  assign T23802 = {T23805, T23803};
  assign T23803 = $signed(T23804) / $signed(22'h100000);
  assign T23804 = $signed(30'h196555b7) * $signed(16'h0);
  assign T23805 = T23803[6'h2d:6'h2d];
  assign T23806 = $signed(T23807) / $signed(22'h100000);
  assign T23807 = $signed(31'h3abee2e5) * $signed(16'h1);
  assign T23808 = T18725[1'h0:1'h0];
  assign T23809 = T23822 ? twiddle4_1_135_real : twiddle4_1_134_real;
  assign twiddle4_1_134_real = T23814 + T23810;
  assign T23810 = {T23813, T23811};
  assign T23811 = $signed(T23812) / $signed(22'h100000);
  assign T23812 = $signed(30'h19937161) * $signed(16'h0);
  assign T23813 = T23811[6'h2d:6'h2d];
  assign T23814 = $signed(T23815) / $signed(22'h100000);
  assign T23815 = $signed(31'h3aaadea5) * $signed(16'h1);
  assign twiddle4_1_135_real = T23820 + T23816;
  assign T23816 = {T23819, T23817};
  assign T23817 = $signed(T23818) / $signed(22'h100000);
  assign T23818 = $signed(30'h19c17d44) * $signed(16'h0);
  assign T23819 = T23817[6'h2d:6'h2d];
  assign T23820 = $signed(T23821) / $signed(22'h100000);
  assign T23821 = $signed(31'h3a96b636) * $signed(16'h1);
  assign T23822 = T18725[1'h0:1'h0];
  assign T23823 = T18725[1'h1:1'h1];
  assign T23824 = T18725[2'h2:2'h2];
  assign T23825 = T23886 ? T23856 : T23826;
  assign T23826 = T23855 ? T23841 : T23827;
  assign T23827 = T23840 ? twiddle4_1_137_real : twiddle4_1_136_real;
  assign twiddle4_1_136_real = T23832 + T23828;
  assign T23828 = {T23831, T23829};
  assign T23829 = $signed(T23830) / $signed(22'h100000);
  assign T23830 = $signed(30'h19ef7943) * $signed(16'h0);
  assign T23831 = T23829[6'h2d:6'h2d];
  assign T23832 = $signed(T23833) / $signed(22'h100000);
  assign T23833 = $signed(31'h3a8269a2) * $signed(16'h1);
  assign twiddle4_1_137_real = T23838 + T23834;
  assign T23834 = {T23837, T23835};
  assign T23835 = $signed(T23836) / $signed(22'h100000);
  assign T23836 = $signed(30'h1a1d6543) * $signed(16'h0);
  assign T23837 = T23835[6'h2d:6'h2d];
  assign T23838 = $signed(T23839) / $signed(22'h100000);
  assign T23839 = $signed(31'h3a6df8f7) * $signed(16'h1);
  assign T23840 = T18725[1'h0:1'h0];
  assign T23841 = T23854 ? twiddle4_1_139_real : twiddle4_1_138_real;
  assign twiddle4_1_138_real = T23846 + T23842;
  assign T23842 = {T23845, T23843};
  assign T23843 = $signed(T23844) / $signed(22'h100000);
  assign T23844 = $signed(30'h1a4b4127) * $signed(16'h0);
  assign T23845 = T23843[6'h2d:6'h2d];
  assign T23846 = $signed(T23847) / $signed(22'h100000);
  assign T23847 = $signed(31'h3a596441) * $signed(16'h1);
  assign twiddle4_1_139_real = T23852 + T23848;
  assign T23848 = {T23851, T23849};
  assign T23849 = $signed(T23850) / $signed(22'h100000);
  assign T23850 = $signed(30'h1a790cd3) * $signed(16'h0);
  assign T23851 = T23849[6'h2d:6'h2d];
  assign T23852 = $signed(T23853) / $signed(22'h100000);
  assign T23853 = $signed(31'h3a44ab8d) * $signed(16'h1);
  assign T23854 = T18725[1'h0:1'h0];
  assign T23855 = T18725[1'h1:1'h1];
  assign T23856 = T23885 ? T23871 : T23857;
  assign T23857 = T23870 ? twiddle4_1_141_real : twiddle4_1_140_real;
  assign twiddle4_1_140_real = T23862 + T23858;
  assign T23858 = {T23861, T23859};
  assign T23859 = $signed(T23860) / $signed(22'h100000);
  assign T23860 = $signed(30'h1aa6c82b) * $signed(16'h0);
  assign T23861 = T23859[6'h2d:6'h2d];
  assign T23862 = $signed(T23863) / $signed(22'h100000);
  assign T23863 = $signed(31'h3a2fcee8) * $signed(16'h1);
  assign twiddle4_1_141_real = T23868 + T23864;
  assign T23864 = {T23867, T23865};
  assign T23865 = $signed(T23866) / $signed(22'h100000);
  assign T23866 = $signed(30'h1ad47312) * $signed(16'h0);
  assign T23867 = T23865[6'h2d:6'h2d];
  assign T23868 = $signed(T23869) / $signed(22'h100000);
  assign T23869 = $signed(31'h3a1ace5e) * $signed(16'h1);
  assign T23870 = T18725[1'h0:1'h0];
  assign T23871 = T23884 ? twiddle4_1_143_real : twiddle4_1_142_real;
  assign twiddle4_1_142_real = T23876 + T23872;
  assign T23872 = {T23875, T23873};
  assign T23873 = $signed(T23874) / $signed(22'h100000);
  assign T23874 = $signed(30'h1b020d6c) * $signed(16'h0);
  assign T23875 = T23873[6'h2d:6'h2d];
  assign T23876 = $signed(T23877) / $signed(22'h100000);
  assign T23877 = $signed(31'h3a05a9fd) * $signed(16'h1);
  assign twiddle4_1_143_real = T23882 + T23878;
  assign T23878 = {T23881, T23879};
  assign T23879 = $signed(T23880) / $signed(22'h100000);
  assign T23880 = $signed(30'h1b2f971d) * $signed(16'h0);
  assign T23881 = T23879[6'h2d:6'h2d];
  assign T23882 = $signed(T23883) / $signed(22'h100000);
  assign T23883 = $signed(31'h39f061d1) * $signed(16'h1);
  assign T23884 = T18725[1'h0:1'h0];
  assign T23885 = T18725[1'h1:1'h1];
  assign T23886 = T18725[2'h2:2'h2];
  assign T23887 = T18725[2'h3:2'h3];
  assign T23888 = T24013 ? T23951 : T23889;
  assign T23889 = T23950 ? T23920 : T23890;
  assign T23890 = T23919 ? T23905 : T23891;
  assign T23891 = T23904 ? twiddle4_1_145_real : twiddle4_1_144_real;
  assign twiddle4_1_144_real = T23896 + T23892;
  assign T23892 = {T23895, T23893};
  assign T23893 = $signed(T23894) / $signed(22'h100000);
  assign T23894 = $signed(30'h1b5d1009) * $signed(16'h0);
  assign T23895 = T23893[6'h2d:6'h2d];
  assign T23896 = $signed(T23897) / $signed(22'h100000);
  assign T23897 = $signed(31'h39daf5e8) * $signed(16'h1);
  assign twiddle4_1_145_real = T23902 + T23898;
  assign T23898 = {T23901, T23899};
  assign T23899 = $signed(T23900) / $signed(22'h100000);
  assign T23900 = $signed(30'h1b8a7814) * $signed(16'h0);
  assign T23901 = T23899[6'h2d:6'h2d];
  assign T23902 = $signed(T23903) / $signed(22'h100000);
  assign T23903 = $signed(31'h39c5664f) * $signed(16'h1);
  assign T23904 = T18725[1'h0:1'h0];
  assign T23905 = T23918 ? twiddle4_1_147_real : twiddle4_1_146_real;
  assign twiddle4_1_146_real = T23910 + T23906;
  assign T23906 = {T23909, T23907};
  assign T23907 = $signed(T23908) / $signed(22'h100000);
  assign T23908 = $signed(30'h1bb7cf23) * $signed(16'h0);
  assign T23909 = T23907[6'h2d:6'h2d];
  assign T23910 = $signed(T23911) / $signed(22'h100000);
  assign T23911 = $signed(31'h39afb313) * $signed(16'h1);
  assign twiddle4_1_147_real = T23916 + T23912;
  assign T23912 = {T23915, T23913};
  assign T23913 = $signed(T23914) / $signed(22'h100000);
  assign T23914 = $signed(30'h1be51517) * $signed(16'h0);
  assign T23915 = T23913[6'h2d:6'h2d];
  assign T23916 = $signed(T23917) / $signed(22'h100000);
  assign T23917 = $signed(31'h3999dc41) * $signed(16'h1);
  assign T23918 = T18725[1'h0:1'h0];
  assign T23919 = T18725[1'h1:1'h1];
  assign T23920 = T23949 ? T23935 : T23921;
  assign T23921 = T23934 ? twiddle4_1_149_real : twiddle4_1_148_real;
  assign twiddle4_1_148_real = T23926 + T23922;
  assign T23922 = {T23925, T23923};
  assign T23923 = $signed(T23924) / $signed(22'h100000);
  assign T23924 = $signed(30'h1c1249d8) * $signed(16'h0);
  assign T23925 = T23923[6'h2d:6'h2d];
  assign T23926 = $signed(T23927) / $signed(22'h100000);
  assign T23927 = $signed(31'h3983e1e7) * $signed(16'h1);
  assign twiddle4_1_149_real = T23932 + T23928;
  assign T23928 = {T23931, T23929};
  assign T23929 = $signed(T23930) / $signed(22'h100000);
  assign T23930 = $signed(30'h1c3f6d47) * $signed(16'h0);
  assign T23931 = T23929[6'h2d:6'h2d];
  assign T23932 = $signed(T23933) / $signed(22'h100000);
  assign T23933 = $signed(31'h396dc414) * $signed(16'h1);
  assign T23934 = T18725[1'h0:1'h0];
  assign T23935 = T23948 ? twiddle4_1_151_real : twiddle4_1_150_real;
  assign twiddle4_1_150_real = T23940 + T23936;
  assign T23936 = {T23939, T23937};
  assign T23937 = $signed(T23938) / $signed(22'h100000);
  assign T23938 = $signed(30'h1c6c7f49) * $signed(16'h0);
  assign T23939 = T23937[6'h2d:6'h2d];
  assign T23940 = $signed(T23941) / $signed(22'h100000);
  assign T23941 = $signed(31'h395782d3) * $signed(16'h1);
  assign twiddle4_1_151_real = T23946 + T23942;
  assign T23942 = {T23945, T23943};
  assign T23943 = $signed(T23944) / $signed(22'h100000);
  assign T23944 = $signed(30'h1c997fc3) * $signed(16'h0);
  assign T23945 = T23943[6'h2d:6'h2d];
  assign T23946 = $signed(T23947) / $signed(22'h100000);
  assign T23947 = $signed(31'h39411e33) * $signed(16'h1);
  assign T23948 = T18725[1'h0:1'h0];
  assign T23949 = T18725[1'h1:1'h1];
  assign T23950 = T18725[2'h2:2'h2];
  assign T23951 = T24012 ? T23982 : T23952;
  assign T23952 = T23981 ? T23967 : T23953;
  assign T23953 = T23966 ? twiddle4_1_153_real : twiddle4_1_152_real;
  assign twiddle4_1_152_real = T23958 + T23954;
  assign T23954 = {T23957, T23955};
  assign T23955 = $signed(T23956) / $signed(22'h100000);
  assign T23956 = $signed(30'h1cc66e99) * $signed(16'h0);
  assign T23957 = T23955[6'h2d:6'h2d];
  assign T23958 = $signed(T23959) / $signed(22'h100000);
  assign T23959 = $signed(31'h392a9642) * $signed(16'h1);
  assign twiddle4_1_153_real = T23964 + T23960;
  assign T23960 = {T23963, T23961};
  assign T23961 = $signed(T23962) / $signed(22'h100000);
  assign T23962 = $signed(30'h1cf34bae) * $signed(16'h0);
  assign T23963 = T23961[6'h2d:6'h2d];
  assign T23964 = $signed(T23965) / $signed(22'h100000);
  assign T23965 = $signed(31'h3913eb0e) * $signed(16'h1);
  assign T23966 = T18725[1'h0:1'h0];
  assign T23967 = T23980 ? twiddle4_1_155_real : twiddle4_1_154_real;
  assign twiddle4_1_154_real = T23972 + T23968;
  assign T23968 = {T23971, T23969};
  assign T23969 = $signed(T23970) / $signed(22'h100000);
  assign T23970 = $signed(30'h1d2016e8) * $signed(16'h0);
  assign T23971 = T23969[6'h2d:6'h2d];
  assign T23972 = $signed(T23973) / $signed(22'h100000);
  assign T23973 = $signed(31'h38fd1ca4) * $signed(16'h1);
  assign twiddle4_1_155_real = T23978 + T23974;
  assign T23974 = {T23977, T23975};
  assign T23975 = $signed(T23976) / $signed(22'h100000);
  assign T23976 = $signed(30'h1d4cd02b) * $signed(16'h0);
  assign T23977 = T23975[6'h2d:6'h2d];
  assign T23978 = $signed(T23979) / $signed(22'h100000);
  assign T23979 = $signed(31'h38e62b13) * $signed(16'h1);
  assign T23980 = T18725[1'h0:1'h0];
  assign T23981 = T18725[1'h1:1'h1];
  assign T23982 = T24011 ? T23997 : T23983;
  assign T23983 = T23996 ? twiddle4_1_157_real : twiddle4_1_156_real;
  assign twiddle4_1_156_real = T23988 + T23984;
  assign T23984 = {T23987, T23985};
  assign T23985 = $signed(T23986) / $signed(22'h100000);
  assign T23986 = $signed(30'h1d79775b) * $signed(16'h0);
  assign T23987 = T23985[6'h2d:6'h2d];
  assign T23988 = $signed(T23989) / $signed(22'h100000);
  assign T23989 = $signed(31'h38cf1669) * $signed(16'h1);
  assign twiddle4_1_157_real = T23994 + T23990;
  assign T23990 = {T23993, T23991};
  assign T23991 = $signed(T23992) / $signed(22'h100000);
  assign T23992 = $signed(30'h1da60c5c) * $signed(16'h0);
  assign T23993 = T23991[6'h2d:6'h2d];
  assign T23994 = $signed(T23995) / $signed(22'h100000);
  assign T23995 = $signed(31'h38b7deb3) * $signed(16'h1);
  assign T23996 = T18725[1'h0:1'h0];
  assign T23997 = T24010 ? twiddle4_1_159_real : twiddle4_1_158_real;
  assign twiddle4_1_158_real = T24002 + T23998;
  assign T23998 = {T24001, T23999};
  assign T23999 = $signed(T24000) / $signed(22'h100000);
  assign T24000 = $signed(30'h1dd28f14) * $signed(16'h0);
  assign T24001 = T23999[6'h2d:6'h2d];
  assign T24002 = $signed(T24003) / $signed(22'h100000);
  assign T24003 = $signed(31'h38a08402) * $signed(16'h1);
  assign twiddle4_1_159_real = T24008 + T24004;
  assign T24004 = {T24007, T24005};
  assign T24005 = $signed(T24006) / $signed(22'h100000);
  assign T24006 = $signed(30'h1dfeff66) * $signed(16'h0);
  assign T24007 = T24005[6'h2d:6'h2d];
  assign T24008 = $signed(T24009) / $signed(22'h100000);
  assign T24009 = $signed(31'h38890662) * $signed(16'h1);
  assign T24010 = T18725[1'h0:1'h0];
  assign T24011 = T18725[1'h1:1'h1];
  assign T24012 = T18725[2'h2:2'h2];
  assign T24013 = T18725[2'h3:2'h3];
  assign T24014 = T18725[3'h4:3'h4];
  assign T24015 = T24226 ? T24132 : T24016;
  assign T24016 = T24131 ? T24079 : T24017;
  assign T24017 = T24078 ? T24048 : T24018;
  assign T24018 = T24047 ? T24033 : T24019;
  assign T24019 = T24032 ? twiddle4_1_161_real : twiddle4_1_160_real;
  assign twiddle4_1_160_real = T24024 + T24020;
  assign T24020 = {T24023, T24021};
  assign T24021 = $signed(T24022) / $signed(22'h100000);
  assign T24022 = $signed(30'h1e2b5d38) * $signed(16'h0);
  assign T24023 = T24021[6'h2d:6'h2d];
  assign T24024 = $signed(T24025) / $signed(22'h100000);
  assign T24025 = $signed(31'h387165e3) * $signed(16'h1);
  assign twiddle4_1_161_real = T24030 + T24026;
  assign T24026 = {T24029, T24027};
  assign T24027 = $signed(T24028) / $signed(22'h100000);
  assign T24028 = $signed(30'h1e57a86d) * $signed(16'h0);
  assign T24029 = T24027[6'h2d:6'h2d];
  assign T24030 = $signed(T24031) / $signed(22'h100000);
  assign T24031 = $signed(31'h3859a292) * $signed(16'h1);
  assign T24032 = T18725[1'h0:1'h0];
  assign T24033 = T24046 ? twiddle4_1_163_real : twiddle4_1_162_real;
  assign twiddle4_1_162_real = T24038 + T24034;
  assign T24034 = {T24037, T24035};
  assign T24035 = $signed(T24036) / $signed(22'h100000);
  assign T24036 = $signed(30'h1e83e0ea) * $signed(16'h0);
  assign T24037 = T24035[6'h2d:6'h2d];
  assign T24038 = $signed(T24039) / $signed(22'h100000);
  assign T24039 = $signed(31'h3841bc7f) * $signed(16'h1);
  assign twiddle4_1_163_real = T24044 + T24040;
  assign T24040 = {T24043, T24041};
  assign T24041 = $signed(T24042) / $signed(22'h100000);
  assign T24042 = $signed(30'h1eb00695) * $signed(16'h0);
  assign T24043 = T24041[6'h2d:6'h2d];
  assign T24044 = $signed(T24045) / $signed(22'h100000);
  assign T24045 = $signed(31'h3829b3b8) * $signed(16'h1);
  assign T24046 = T18725[1'h0:1'h0];
  assign T24047 = T18725[1'h1:1'h1];
  assign T24048 = T24077 ? T24063 : T24049;
  assign T24049 = T24062 ? twiddle4_1_165_real : twiddle4_1_164_real;
  assign twiddle4_1_164_real = T24054 + T24050;
  assign T24050 = {T24053, T24051};
  assign T24051 = $signed(T24052) / $signed(22'h100000);
  assign T24052 = $signed(30'h1edc1952) * $signed(16'h0);
  assign T24053 = T24051[6'h2d:6'h2d];
  assign T24054 = $signed(T24055) / $signed(22'h100000);
  assign T24055 = $signed(31'h3811884c) * $signed(16'h1);
  assign twiddle4_1_165_real = T24060 + T24056;
  assign T24056 = {T24059, T24057};
  assign T24057 = $signed(T24058) / $signed(22'h100000);
  assign T24058 = $signed(30'h1f081906) * $signed(16'h0);
  assign T24059 = T24057[6'h2d:6'h2d];
  assign T24060 = $signed(T24061) / $signed(22'h100000);
  assign T24061 = $signed(31'h37f93a4b) * $signed(16'h1);
  assign T24062 = T18725[1'h0:1'h0];
  assign T24063 = T24076 ? twiddle4_1_167_real : twiddle4_1_166_real;
  assign twiddle4_1_166_real = T24068 + T24064;
  assign T24064 = {T24067, T24065};
  assign T24065 = $signed(T24066) / $signed(22'h100000);
  assign T24066 = $signed(30'h1f340596) * $signed(16'h0);
  assign T24067 = T24065[6'h2d:6'h2d];
  assign T24068 = $signed(T24069) / $signed(22'h100000);
  assign T24069 = $signed(31'h37e0c9c2) * $signed(16'h1);
  assign twiddle4_1_167_real = T24074 + T24070;
  assign T24070 = {T24073, T24071};
  assign T24071 = $signed(T24072) / $signed(22'h100000);
  assign T24072 = $signed(30'h1f5fdee6) * $signed(16'h0);
  assign T24073 = T24071[6'h2d:6'h2d];
  assign T24074 = $signed(T24075) / $signed(22'h100000);
  assign T24075 = $signed(31'h37c836c2) * $signed(16'h1);
  assign T24076 = T18725[1'h0:1'h0];
  assign T24077 = T18725[1'h1:1'h1];
  assign T24078 = T18725[2'h2:2'h2];
  assign T24079 = T24130 ? T24108 : T24080;
  assign T24080 = T24107 ? T24095 : T24081;
  assign T24081 = T24094 ? twiddle4_1_169_real : twiddle4_1_168_real;
  assign twiddle4_1_168_real = T24086 + T24082;
  assign T24082 = {T24085, T24083};
  assign T24083 = $signed(T24084) / $signed(22'h100000);
  assign T24084 = $signed(30'h1f8ba4db) * $signed(16'h0);
  assign T24085 = T24083[6'h2d:6'h2d];
  assign T24086 = $signed(T24087) / $signed(22'h100000);
  assign T24087 = $signed(31'h37af8158) * $signed(16'h1);
  assign twiddle4_1_169_real = T24092 + T24088;
  assign T24088 = {T24091, T24089};
  assign T24089 = $signed(T24090) / $signed(22'h100000);
  assign T24090 = $signed(30'h1fb7575c) * $signed(16'h0);
  assign T24091 = T24089[6'h2d:6'h2d];
  assign T24092 = $signed(T24093) / $signed(22'h100000);
  assign T24093 = $signed(31'h3796a996) * $signed(16'h1);
  assign T24094 = T18725[1'h0:1'h0];
  assign T24095 = T24106 ? twiddle4_1_171_real : twiddle4_1_170_real;
  assign twiddle4_1_170_real = T24100 + T24096;
  assign T24096 = {T24099, T24097};
  assign T24097 = $signed(T24098) / $signed(22'h100000);
  assign T24098 = $signed(30'h1fe2f64b) * $signed(16'h0);
  assign T24099 = T24097[6'h2d:6'h2d];
  assign T24100 = $signed(T24101) / $signed(22'h100000);
  assign T24101 = $signed(31'h377daf89) * $signed(16'h1);
  assign twiddle4_1_171_real = T24104 + T24102;
  assign T24102 = $signed(T24103) / $signed(22'h100000);
  assign T24103 = $signed(31'h200e8190) * $signed(16'h0);
  assign T24104 = $signed(T24105) / $signed(22'h100000);
  assign T24105 = $signed(31'h37649341) * $signed(16'h1);
  assign T24106 = T18725[1'h0:1'h0];
  assign T24107 = T18725[1'h1:1'h1];
  assign T24108 = T24129 ? T24119 : T24109;
  assign T24109 = T24118 ? twiddle4_1_173_real : twiddle4_1_172_real;
  assign twiddle4_1_172_real = T24112 + T24110;
  assign T24110 = $signed(T24111) / $signed(22'h100000);
  assign T24111 = $signed(31'h2039f90e) * $signed(16'h0);
  assign T24112 = $signed(T24113) / $signed(22'h100000);
  assign T24113 = $signed(31'h374b54ce) * $signed(16'h1);
  assign twiddle4_1_173_real = T24116 + T24114;
  assign T24114 = $signed(T24115) / $signed(22'h100000);
  assign T24115 = $signed(31'h20655cab) * $signed(16'h0);
  assign T24116 = $signed(T24117) / $signed(22'h100000);
  assign T24117 = $signed(31'h3731f43f) * $signed(16'h1);
  assign T24118 = T18725[1'h0:1'h0];
  assign T24119 = T24128 ? twiddle4_1_175_real : twiddle4_1_174_real;
  assign twiddle4_1_174_real = T24122 + T24120;
  assign T24120 = $signed(T24121) / $signed(22'h100000);
  assign T24121 = $signed(31'h2090ac4d) * $signed(16'h0);
  assign T24122 = $signed(T24123) / $signed(22'h100000);
  assign T24123 = $signed(31'h371871a4) * $signed(16'h1);
  assign twiddle4_1_175_real = T24126 + T24124;
  assign T24124 = $signed(T24125) / $signed(22'h100000);
  assign T24125 = $signed(31'h20bbe7d8) * $signed(16'h0);
  assign T24126 = $signed(T24127) / $signed(22'h100000);
  assign T24127 = $signed(31'h36fecd0d) * $signed(16'h1);
  assign T24128 = T18725[1'h0:1'h0];
  assign T24129 = T18725[1'h1:1'h1];
  assign T24130 = T18725[2'h2:2'h2];
  assign T24131 = T18725[2'h3:2'h3];
  assign T24132 = T24225 ? T24179 : T24133;
  assign T24133 = T24178 ? T24156 : T24134;
  assign T24134 = T24155 ? T24145 : T24135;
  assign T24135 = T24144 ? twiddle4_1_177_real : twiddle4_1_176_real;
  assign twiddle4_1_176_real = T24138 + T24136;
  assign T24136 = $signed(T24137) / $signed(22'h100000);
  assign T24137 = $signed(31'h20e70f32) * $signed(16'h0);
  assign T24138 = $signed(T24139) / $signed(22'h100000);
  assign T24139 = $signed(31'h36e5068a) * $signed(16'h1);
  assign twiddle4_1_177_real = T24142 + T24140;
  assign T24140 = $signed(T24141) / $signed(22'h100000);
  assign T24141 = $signed(31'h21122240) * $signed(16'h0);
  assign T24142 = $signed(T24143) / $signed(22'h100000);
  assign T24143 = $signed(31'h36cb1e29) * $signed(16'h1);
  assign T24144 = T18725[1'h0:1'h0];
  assign T24145 = T24154 ? twiddle4_1_179_real : twiddle4_1_178_real;
  assign twiddle4_1_178_real = T24148 + T24146;
  assign T24146 = $signed(T24147) / $signed(22'h100000);
  assign T24147 = $signed(31'h213d20e8) * $signed(16'h0);
  assign T24148 = $signed(T24149) / $signed(22'h100000);
  assign T24149 = $signed(31'h36b113fd) * $signed(16'h1);
  assign twiddle4_1_179_real = T24152 + T24150;
  assign T24150 = $signed(T24151) / $signed(22'h100000);
  assign T24151 = $signed(31'h21680b0f) * $signed(16'h0);
  assign T24152 = $signed(T24153) / $signed(22'h100000);
  assign T24153 = $signed(31'h3696e813) * $signed(16'h1);
  assign T24154 = T18725[1'h0:1'h0];
  assign T24155 = T18725[1'h1:1'h1];
  assign T24156 = T24177 ? T24167 : T24157;
  assign T24157 = T24166 ? twiddle4_1_181_real : twiddle4_1_180_real;
  assign twiddle4_1_180_real = T24160 + T24158;
  assign T24158 = $signed(T24159) / $signed(22'h100000);
  assign T24159 = $signed(31'h2192e09a) * $signed(16'h0);
  assign T24160 = $signed(T24161) / $signed(22'h100000);
  assign T24161 = $signed(31'h367c9a7d) * $signed(16'h1);
  assign twiddle4_1_181_real = T24164 + T24162;
  assign T24162 = $signed(T24163) / $signed(22'h100000);
  assign T24163 = $signed(31'h21bda170) * $signed(16'h0);
  assign T24164 = $signed(T24165) / $signed(22'h100000);
  assign T24165 = $signed(31'h36622b4b) * $signed(16'h1);
  assign T24166 = T18725[1'h0:1'h0];
  assign T24167 = T24176 ? twiddle4_1_183_real : twiddle4_1_182_real;
  assign twiddle4_1_182_real = T24170 + T24168;
  assign T24168 = $signed(T24169) / $signed(22'h100000);
  assign T24169 = $signed(31'h21e84d76) * $signed(16'h0);
  assign T24170 = $signed(T24171) / $signed(22'h100000);
  assign T24171 = $signed(31'h36479a8e) * $signed(16'h1);
  assign twiddle4_1_183_real = T24174 + T24172;
  assign T24172 = $signed(T24173) / $signed(22'h100000);
  assign T24173 = $signed(31'h2212e491) * $signed(16'h0);
  assign T24174 = $signed(T24175) / $signed(22'h100000);
  assign T24175 = $signed(31'h362ce854) * $signed(16'h1);
  assign T24176 = T18725[1'h0:1'h0];
  assign T24177 = T18725[1'h1:1'h1];
  assign T24178 = T18725[2'h2:2'h2];
  assign T24179 = T24224 ? T24202 : T24180;
  assign T24180 = T24201 ? T24191 : T24181;
  assign T24181 = T24190 ? twiddle4_1_185_real : twiddle4_1_184_real;
  assign twiddle4_1_184_real = T24184 + T24182;
  assign T24182 = $signed(T24183) / $signed(22'h100000);
  assign T24183 = $signed(31'h223d66a8) * $signed(16'h0);
  assign T24184 = $signed(T24185) / $signed(22'h100000);
  assign T24185 = $signed(31'h361214b0) * $signed(16'h1);
  assign twiddle4_1_185_real = T24188 + T24186;
  assign T24186 = $signed(T24187) / $signed(22'h100000);
  assign T24187 = $signed(31'h2267d39f) * $signed(16'h0);
  assign T24188 = $signed(T24189) / $signed(22'h100000);
  assign T24189 = $signed(31'h35f71fb1) * $signed(16'h1);
  assign T24190 = T18725[1'h0:1'h0];
  assign T24191 = T24200 ? twiddle4_1_187_real : twiddle4_1_186_real;
  assign twiddle4_1_186_real = T24194 + T24192;
  assign T24192 = $signed(T24193) / $signed(22'h100000);
  assign T24193 = $signed(31'h22922b5e) * $signed(16'h0);
  assign T24194 = $signed(T24195) / $signed(22'h100000);
  assign T24195 = $signed(31'h35dc0968) * $signed(16'h1);
  assign twiddle4_1_187_real = T24198 + T24196;
  assign T24196 = $signed(T24197) / $signed(22'h100000);
  assign T24197 = $signed(31'h22bc6dc9) * $signed(16'h0);
  assign T24198 = $signed(T24199) / $signed(22'h100000);
  assign T24199 = $signed(31'h35c0d1e6) * $signed(16'h1);
  assign T24200 = T18725[1'h0:1'h0];
  assign T24201 = T18725[1'h1:1'h1];
  assign T24202 = T24223 ? T24213 : T24203;
  assign T24203 = T24212 ? twiddle4_1_189_real : twiddle4_1_188_real;
  assign twiddle4_1_188_real = T24206 + T24204;
  assign T24204 = $signed(T24205) / $signed(22'h100000);
  assign T24205 = $signed(31'h22e69ac7) * $signed(16'h0);
  assign T24206 = $signed(T24207) / $signed(22'h100000);
  assign T24207 = $signed(31'h35a5793c) * $signed(16'h1);
  assign twiddle4_1_189_real = T24210 + T24208;
  assign T24208 = $signed(T24209) / $signed(22'h100000);
  assign T24209 = $signed(31'h2310b23e) * $signed(16'h0);
  assign T24210 = $signed(T24211) / $signed(22'h100000);
  assign T24211 = $signed(31'h3589ff7a) * $signed(16'h1);
  assign T24212 = T18725[1'h0:1'h0];
  assign T24213 = T24222 ? twiddle4_1_191_real : twiddle4_1_190_real;
  assign twiddle4_1_190_real = T24216 + T24214;
  assign T24214 = $signed(T24215) / $signed(22'h100000);
  assign T24215 = $signed(31'h233ab413) * $signed(16'h0);
  assign T24216 = $signed(T24217) / $signed(22'h100000);
  assign T24217 = $signed(31'h356e64b2) * $signed(16'h1);
  assign twiddle4_1_191_real = T24220 + T24218;
  assign T24218 = $signed(T24219) / $signed(22'h100000);
  assign T24219 = $signed(31'h2364a02e) * $signed(16'h0);
  assign T24220 = $signed(T24221) / $signed(22'h100000);
  assign T24221 = $signed(31'h3552a8f4) * $signed(16'h1);
  assign T24222 = T18725[1'h0:1'h0];
  assign T24223 = T18725[1'h1:1'h1];
  assign T24224 = T18725[2'h2:2'h2];
  assign T24225 = T18725[2'h3:2'h3];
  assign T24226 = T18725[3'h4:3'h4];
  assign T24227 = T18725[3'h5:3'h5];
  assign T24228 = T24609 ? T24419 : T24229;
  assign T24229 = T24418 ? T24324 : T24230;
  assign T24230 = T24323 ? T24277 : T24231;
  assign T24231 = T24276 ? T24254 : T24232;
  assign T24232 = T24253 ? T24243 : T24233;
  assign T24233 = T24242 ? twiddle4_1_193_real : twiddle4_1_192_real;
  assign twiddle4_1_192_real = T24236 + T24234;
  assign T24234 = $signed(T24235) / $signed(22'h100000);
  assign T24235 = $signed(31'h238e7673) * $signed(16'h0);
  assign T24236 = $signed(T24237) / $signed(22'h100000);
  assign T24237 = $signed(31'h3536cc52) * $signed(16'h1);
  assign twiddle4_1_193_real = T24240 + T24238;
  assign T24238 = $signed(T24239) / $signed(22'h100000);
  assign T24239 = $signed(31'h23b836c9) * $signed(16'h0);
  assign T24240 = $signed(T24241) / $signed(22'h100000);
  assign T24241 = $signed(31'h351acedc) * $signed(16'h1);
  assign T24242 = T18725[1'h0:1'h0];
  assign T24243 = T24252 ? twiddle4_1_195_real : twiddle4_1_194_real;
  assign twiddle4_1_194_real = T24246 + T24244;
  assign T24244 = $signed(T24245) / $signed(22'h100000);
  assign T24245 = $signed(31'h23e1e117) * $signed(16'h0);
  assign T24246 = $signed(T24247) / $signed(22'h100000);
  assign T24247 = $signed(31'h34feb0a5) * $signed(16'h1);
  assign twiddle4_1_195_real = T24250 + T24248;
  assign T24248 = $signed(T24249) / $signed(22'h100000);
  assign T24249 = $signed(31'h240b7542) * $signed(16'h0);
  assign T24250 = $signed(T24251) / $signed(22'h100000);
  assign T24251 = $signed(31'h34e271bd) * $signed(16'h1);
  assign T24252 = T18725[1'h0:1'h0];
  assign T24253 = T18725[1'h1:1'h1];
  assign T24254 = T24275 ? T24265 : T24255;
  assign T24255 = T24264 ? twiddle4_1_197_real : twiddle4_1_196_real;
  assign twiddle4_1_196_real = T24258 + T24256;
  assign T24256 = $signed(T24257) / $signed(22'h100000);
  assign T24257 = $signed(31'h2434f332) * $signed(16'h0);
  assign T24258 = $signed(T24259) / $signed(22'h100000);
  assign T24259 = $signed(31'h34c61236) * $signed(16'h1);
  assign twiddle4_1_197_real = T24262 + T24260;
  assign T24260 = $signed(T24261) / $signed(22'h100000);
  assign T24261 = $signed(31'h245e5acc) * $signed(16'h0);
  assign T24262 = $signed(T24263) / $signed(22'h100000);
  assign T24263 = $signed(31'h34a99221) * $signed(16'h1);
  assign T24264 = T18725[1'h0:1'h0];
  assign T24265 = T24274 ? twiddle4_1_199_real : twiddle4_1_198_real;
  assign twiddle4_1_198_real = T24268 + T24266;
  assign T24266 = $signed(T24267) / $signed(22'h100000);
  assign T24267 = $signed(31'h2487abf7) * $signed(16'h0);
  assign T24268 = $signed(T24269) / $signed(22'h100000);
  assign T24269 = $signed(31'h348cf190) * $signed(16'h1);
  assign twiddle4_1_199_real = T24272 + T24270;
  assign T24270 = $signed(T24271) / $signed(22'h100000);
  assign T24271 = $signed(31'h24b0e699) * $signed(16'h0);
  assign T24272 = $signed(T24273) / $signed(22'h100000);
  assign T24273 = $signed(31'h34703094) * $signed(16'h1);
  assign T24274 = T18725[1'h0:1'h0];
  assign T24275 = T18725[1'h1:1'h1];
  assign T24276 = T18725[2'h2:2'h2];
  assign T24277 = T24322 ? T24300 : T24278;
  assign T24278 = T24299 ? T24289 : T24279;
  assign T24279 = T24288 ? twiddle4_1_201_real : twiddle4_1_200_real;
  assign twiddle4_1_200_real = T24282 + T24280;
  assign T24280 = $signed(T24281) / $signed(22'h100000);
  assign T24281 = $signed(31'h24da0a99) * $signed(16'h0);
  assign T24282 = $signed(T24283) / $signed(22'h100000);
  assign T24283 = $signed(31'h34534f40) * $signed(16'h1);
  assign twiddle4_1_201_real = T24286 + T24284;
  assign T24284 = $signed(T24285) / $signed(22'h100000);
  assign T24285 = $signed(31'h250317de) * $signed(16'h0);
  assign T24286 = $signed(T24287) / $signed(22'h100000);
  assign T24287 = $signed(31'h34364da5) * $signed(16'h1);
  assign T24288 = T18725[1'h0:1'h0];
  assign T24289 = T24298 ? twiddle4_1_203_real : twiddle4_1_202_real;
  assign twiddle4_1_202_real = T24292 + T24290;
  assign T24290 = $signed(T24291) / $signed(22'h100000);
  assign T24291 = $signed(31'h252c0e4e) * $signed(16'h0);
  assign T24292 = $signed(T24293) / $signed(22'h100000);
  assign T24293 = $signed(31'h34192bd5) * $signed(16'h1);
  assign twiddle4_1_203_real = T24296 + T24294;
  assign T24294 = $signed(T24295) / $signed(22'h100000);
  assign T24295 = $signed(31'h2554edd0) * $signed(16'h0);
  assign T24296 = $signed(T24297) / $signed(22'h100000);
  assign T24297 = $signed(31'h33fbe9e2) * $signed(16'h1);
  assign T24298 = T18725[1'h0:1'h0];
  assign T24299 = T18725[1'h1:1'h1];
  assign T24300 = T24321 ? T24311 : T24301;
  assign T24301 = T24310 ? twiddle4_1_205_real : twiddle4_1_204_real;
  assign twiddle4_1_204_real = T24304 + T24302;
  assign T24302 = $signed(T24303) / $signed(22'h100000);
  assign T24303 = $signed(31'h257db64b) * $signed(16'h0);
  assign T24304 = $signed(T24305) / $signed(22'h100000);
  assign T24305 = $signed(31'h33de87de) * $signed(16'h1);
  assign twiddle4_1_205_real = T24308 + T24306;
  assign T24306 = $signed(T24307) / $signed(22'h100000);
  assign T24307 = $signed(31'h25a667a6) * $signed(16'h0);
  assign T24308 = $signed(T24309) / $signed(22'h100000);
  assign T24309 = $signed(31'h33c105db) * $signed(16'h1);
  assign T24310 = T18725[1'h0:1'h0];
  assign T24311 = T24320 ? twiddle4_1_207_real : twiddle4_1_206_real;
  assign twiddle4_1_206_real = T24314 + T24312;
  assign T24312 = $signed(T24313) / $signed(22'h100000);
  assign T24313 = $signed(31'h25cf01c7) * $signed(16'h0);
  assign T24314 = $signed(T24315) / $signed(22'h100000);
  assign T24315 = $signed(31'h33a363eb) * $signed(16'h1);
  assign twiddle4_1_207_real = T24318 + T24316;
  assign T24316 = $signed(T24317) / $signed(22'h100000);
  assign T24317 = $signed(31'h25f78496) * $signed(16'h0);
  assign T24318 = $signed(T24319) / $signed(22'h100000);
  assign T24319 = $signed(31'h3385a221) * $signed(16'h1);
  assign T24320 = T18725[1'h0:1'h0];
  assign T24321 = T18725[1'h1:1'h1];
  assign T24322 = T18725[2'h2:2'h2];
  assign T24323 = T18725[2'h3:2'h3];
  assign T24324 = T24417 ? T24371 : T24325;
  assign T24325 = T24370 ? T24348 : T24326;
  assign T24326 = T24347 ? T24337 : T24327;
  assign T24327 = T24336 ? twiddle4_1_209_real : twiddle4_1_208_real;
  assign twiddle4_1_208_real = T24330 + T24328;
  assign T24328 = $signed(T24329) / $signed(22'h100000);
  assign T24329 = $signed(31'h261feff9) * $signed(16'h0);
  assign T24330 = $signed(T24331) / $signed(22'h100000);
  assign T24331 = $signed(31'h3367c08f) * $signed(16'h1);
  assign twiddle4_1_209_real = T24334 + T24332;
  assign T24332 = $signed(T24333) / $signed(22'h100000);
  assign T24333 = $signed(31'h264843d8) * $signed(16'h0);
  assign T24334 = $signed(T24335) / $signed(22'h100000);
  assign T24335 = $signed(31'h3349bf48) * $signed(16'h1);
  assign T24336 = T18725[1'h0:1'h0];
  assign T24337 = T24346 ? twiddle4_1_211_real : twiddle4_1_210_real;
  assign twiddle4_1_210_real = T24340 + T24338;
  assign T24338 = $signed(T24339) / $signed(22'h100000);
  assign T24339 = $signed(31'h2670801a) * $signed(16'h0);
  assign T24340 = $signed(T24341) / $signed(22'h100000);
  assign T24341 = $signed(31'h332b9e5d) * $signed(16'h1);
  assign twiddle4_1_211_real = T24344 + T24342;
  assign T24342 = $signed(T24343) / $signed(22'h100000);
  assign T24343 = $signed(31'h2698a4a5) * $signed(16'h0);
  assign T24344 = $signed(T24345) / $signed(22'h100000);
  assign T24345 = $signed(31'h330d5de2) * $signed(16'h1);
  assign T24346 = T18725[1'h0:1'h0];
  assign T24347 = T18725[1'h1:1'h1];
  assign T24348 = T24369 ? T24359 : T24349;
  assign T24349 = T24358 ? twiddle4_1_213_real : twiddle4_1_212_real;
  assign twiddle4_1_212_real = T24352 + T24350;
  assign T24350 = $signed(T24351) / $signed(22'h100000);
  assign T24351 = $signed(31'h26c0b162) * $signed(16'h0);
  assign T24352 = $signed(T24353) / $signed(22'h100000);
  assign T24353 = $signed(31'h32eefde9) * $signed(16'h1);
  assign twiddle4_1_213_real = T24356 + T24354;
  assign T24354 = $signed(T24355) / $signed(22'h100000);
  assign T24355 = $signed(31'h26e8a637) * $signed(16'h0);
  assign T24356 = $signed(T24357) / $signed(22'h100000);
  assign T24357 = $signed(31'h32d07e85) * $signed(16'h1);
  assign T24358 = T18725[1'h0:1'h0];
  assign T24359 = T24368 ? twiddle4_1_215_real : twiddle4_1_214_real;
  assign twiddle4_1_214_real = T24362 + T24360;
  assign T24360 = $signed(T24361) / $signed(22'h100000);
  assign T24361 = $signed(31'h2710830b) * $signed(16'h0);
  assign T24362 = $signed(T24363) / $signed(22'h100000);
  assign T24363 = $signed(31'h32b1dfc9) * $signed(16'h1);
  assign twiddle4_1_215_real = T24366 + T24364;
  assign T24364 = $signed(T24365) / $signed(22'h100000);
  assign T24365 = $signed(31'h273847c7) * $signed(16'h0);
  assign T24366 = $signed(T24367) / $signed(22'h100000);
  assign T24367 = $signed(31'h329321c7) * $signed(16'h1);
  assign T24368 = T18725[1'h0:1'h0];
  assign T24369 = T18725[1'h1:1'h1];
  assign T24370 = T18725[2'h2:2'h2];
  assign T24371 = T24416 ? T24394 : T24372;
  assign T24372 = T24393 ? T24383 : T24373;
  assign T24373 = T24382 ? twiddle4_1_217_real : twiddle4_1_216_real;
  assign twiddle4_1_216_real = T24376 + T24374;
  assign T24374 = $signed(T24375) / $signed(22'h100000);
  assign T24375 = $signed(31'h275ff452) * $signed(16'h0);
  assign T24376 = $signed(T24377) / $signed(22'h100000);
  assign T24377 = $signed(31'h32744493) * $signed(16'h1);
  assign twiddle4_1_217_real = T24380 + T24378;
  assign T24378 = $signed(T24379) / $signed(22'h100000);
  assign T24379 = $signed(31'h27878893) * $signed(16'h0);
  assign T24380 = $signed(T24381) / $signed(22'h100000);
  assign T24381 = $signed(31'h3255483f) * $signed(16'h1);
  assign T24382 = T18725[1'h0:1'h0];
  assign T24383 = T24392 ? twiddle4_1_219_real : twiddle4_1_218_real;
  assign twiddle4_1_218_real = T24386 + T24384;
  assign T24384 = $signed(T24385) / $signed(22'h100000);
  assign T24385 = $signed(31'h27af0471) * $signed(16'h0);
  assign T24386 = $signed(T24387) / $signed(22'h100000);
  assign T24387 = $signed(31'h32362cdf) * $signed(16'h1);
  assign twiddle4_1_219_real = T24390 + T24388;
  assign T24388 = $signed(T24389) / $signed(22'h100000);
  assign T24389 = $signed(31'h27d667d5) * $signed(16'h0);
  assign T24390 = $signed(T24391) / $signed(22'h100000);
  assign T24391 = $signed(31'h3216f286) * $signed(16'h1);
  assign T24392 = T18725[1'h0:1'h0];
  assign T24393 = T18725[1'h1:1'h1];
  assign T24394 = T24415 ? T24405 : T24395;
  assign T24395 = T24404 ? twiddle4_1_221_real : twiddle4_1_220_real;
  assign twiddle4_1_220_real = T24398 + T24396;
  assign T24396 = $signed(T24397) / $signed(22'h100000);
  assign T24397 = $signed(31'h27fdb2a6) * $signed(16'h0);
  assign T24398 = $signed(T24399) / $signed(22'h100000);
  assign T24399 = $signed(31'h31f79947) * $signed(16'h1);
  assign twiddle4_1_221_real = T24402 + T24400;
  assign T24400 = $signed(T24401) / $signed(22'h100000);
  assign T24401 = $signed(31'h2824e4cc) * $signed(16'h0);
  assign T24402 = $signed(T24403) / $signed(22'h100000);
  assign T24403 = $signed(31'h31d82136) * $signed(16'h1);
  assign T24404 = T18725[1'h0:1'h0];
  assign T24405 = T24414 ? twiddle4_1_223_real : twiddle4_1_222_real;
  assign twiddle4_1_222_real = T24408 + T24406;
  assign T24406 = $signed(T24407) / $signed(22'h100000);
  assign T24407 = $signed(31'h284bfe2f) * $signed(16'h0);
  assign T24408 = $signed(T24409) / $signed(22'h100000);
  assign T24409 = $signed(31'h31b88a66) * $signed(16'h1);
  assign twiddle4_1_223_real = T24412 + T24410;
  assign T24410 = $signed(T24411) / $signed(22'h100000);
  assign T24411 = $signed(31'h2872feb6) * $signed(16'h0);
  assign T24412 = $signed(T24413) / $signed(22'h100000);
  assign T24413 = $signed(31'h3198d4ea) * $signed(16'h1);
  assign T24414 = T18725[1'h0:1'h0];
  assign T24415 = T18725[1'h1:1'h1];
  assign T24416 = T18725[2'h2:2'h2];
  assign T24417 = T18725[2'h3:2'h3];
  assign T24418 = T18725[3'h4:3'h4];
  assign T24419 = T24608 ? T24514 : T24420;
  assign T24420 = T24513 ? T24467 : T24421;
  assign T24421 = T24466 ? T24444 : T24422;
  assign T24422 = T24443 ? T24433 : T24423;
  assign T24423 = T24432 ? twiddle4_1_225_real : twiddle4_1_224_real;
  assign twiddle4_1_224_real = T24426 + T24424;
  assign T24424 = $signed(T24425) / $signed(22'h100000);
  assign T24425 = $signed(31'h2899e64a) * $signed(16'h0);
  assign T24426 = $signed(T24427) / $signed(22'h100000);
  assign T24427 = $signed(31'h317900d6) * $signed(16'h1);
  assign twiddle4_1_225_real = T24430 + T24428;
  assign T24428 = $signed(T24429) / $signed(22'h100000);
  assign T24429 = $signed(31'h28c0b4d2) * $signed(16'h0);
  assign T24430 = $signed(T24431) / $signed(22'h100000);
  assign T24431 = $signed(31'h31590e3d) * $signed(16'h1);
  assign T24432 = T18725[1'h0:1'h0];
  assign T24433 = T24442 ? twiddle4_1_227_real : twiddle4_1_226_real;
  assign twiddle4_1_226_real = T24436 + T24434;
  assign T24434 = $signed(T24435) / $signed(22'h100000);
  assign T24435 = $signed(31'h28e76a37) * $signed(16'h0);
  assign T24436 = $signed(T24437) / $signed(22'h100000);
  assign T24437 = $signed(31'h3138fd34) * $signed(16'h1);
  assign twiddle4_1_227_real = T24440 + T24438;
  assign T24438 = $signed(T24439) / $signed(22'h100000);
  assign T24439 = $signed(31'h290e0660) * $signed(16'h0);
  assign T24440 = $signed(T24441) / $signed(22'h100000);
  assign T24441 = $signed(31'h3118cdce) * $signed(16'h1);
  assign T24442 = T18725[1'h0:1'h0];
  assign T24443 = T18725[1'h1:1'h1];
  assign T24444 = T24465 ? T24455 : T24445;
  assign T24445 = T24454 ? twiddle4_1_229_real : twiddle4_1_228_real;
  assign twiddle4_1_228_real = T24448 + T24446;
  assign T24446 = $signed(T24447) / $signed(22'h100000);
  assign T24447 = $signed(31'h29348937) * $signed(16'h0);
  assign T24448 = $signed(T24449) / $signed(22'h100000);
  assign T24449 = $signed(31'h30f8801f) * $signed(16'h1);
  assign twiddle4_1_229_real = T24452 + T24450;
  assign T24450 = $signed(T24451) / $signed(22'h100000);
  assign T24451 = $signed(31'h295af2a2) * $signed(16'h0);
  assign T24452 = $signed(T24453) / $signed(22'h100000);
  assign T24453 = $signed(31'h30d8143b) * $signed(16'h1);
  assign T24454 = T18725[1'h0:1'h0];
  assign T24455 = T24464 ? twiddle4_1_231_real : twiddle4_1_230_real;
  assign twiddle4_1_230_real = T24458 + T24456;
  assign T24456 = $signed(T24457) / $signed(22'h100000);
  assign T24457 = $signed(31'h2981428b) * $signed(16'h0);
  assign T24458 = $signed(T24459) / $signed(22'h100000);
  assign T24459 = $signed(31'h30b78a35) * $signed(16'h1);
  assign twiddle4_1_231_real = T24462 + T24460;
  assign T24460 = $signed(T24461) / $signed(22'h100000);
  assign T24461 = $signed(31'h29a778da) * $signed(16'h0);
  assign T24462 = $signed(T24463) / $signed(22'h100000);
  assign T24463 = $signed(31'h3096e223) * $signed(16'h1);
  assign T24464 = T18725[1'h0:1'h0];
  assign T24465 = T18725[1'h1:1'h1];
  assign T24466 = T18725[2'h2:2'h2];
  assign T24467 = T24512 ? T24490 : T24468;
  assign T24468 = T24489 ? T24479 : T24469;
  assign T24469 = T24478 ? twiddle4_1_233_real : twiddle4_1_232_real;
  assign twiddle4_1_232_real = T24472 + T24470;
  assign T24470 = $signed(T24471) / $signed(22'h100000);
  assign T24471 = $signed(31'h29cd9577) * $signed(16'h0);
  assign T24472 = $signed(T24473) / $signed(22'h100000);
  assign T24473 = $signed(31'h30761c17) * $signed(16'h1);
  assign twiddle4_1_233_real = T24476 + T24474;
  assign T24474 = $signed(T24475) / $signed(22'h100000);
  assign T24475 = $signed(31'h29f3984b) * $signed(16'h0);
  assign T24476 = $signed(T24477) / $signed(22'h100000);
  assign T24477 = $signed(31'h30553827) * $signed(16'h1);
  assign T24478 = T18725[1'h0:1'h0];
  assign T24479 = T24488 ? twiddle4_1_235_real : twiddle4_1_234_real;
  assign twiddle4_1_234_real = T24482 + T24480;
  assign T24480 = $signed(T24481) / $signed(22'h100000);
  assign T24481 = $signed(31'h2a19813e) * $signed(16'h0);
  assign T24482 = $signed(T24483) / $signed(22'h100000);
  assign T24483 = $signed(31'h30343667) * $signed(16'h1);
  assign twiddle4_1_235_real = T24486 + T24484;
  assign T24484 = $signed(T24485) / $signed(22'h100000);
  assign T24485 = $signed(31'h2a3f5039) * $signed(16'h0);
  assign T24486 = $signed(T24487) / $signed(22'h100000);
  assign T24487 = $signed(31'h301316ea) * $signed(16'h1);
  assign T24488 = T18725[1'h0:1'h0];
  assign T24489 = T18725[1'h1:1'h1];
  assign T24490 = T24511 ? T24501 : T24491;
  assign T24491 = T24500 ? twiddle4_1_237_real : twiddle4_1_236_real;
  assign twiddle4_1_236_real = T24494 + T24492;
  assign T24492 = $signed(T24493) / $signed(22'h100000);
  assign T24493 = $signed(31'h2a650525) * $signed(16'h0);
  assign T24494 = $signed(T24495) / $signed(22'h100000);
  assign T24495 = $signed(31'h2ff1d9c6) * $signed(16'h1);
  assign twiddle4_1_237_real = T24498 + T24496;
  assign T24496 = $signed(T24497) / $signed(22'h100000);
  assign T24497 = $signed(31'h2a8a9fea) * $signed(16'h0);
  assign T24498 = $signed(T24499) / $signed(22'h100000);
  assign T24499 = $signed(31'h2fd07f0f) * $signed(16'h1);
  assign T24500 = T18725[1'h0:1'h0];
  assign T24501 = T24510 ? twiddle4_1_239_real : twiddle4_1_238_real;
  assign twiddle4_1_238_real = T24504 + T24502;
  assign T24502 = $signed(T24503) / $signed(22'h100000);
  assign T24503 = $signed(31'h2ab02071) * $signed(16'h0);
  assign T24504 = $signed(T24505) / $signed(22'h100000);
  assign T24505 = $signed(31'h2faf06d9) * $signed(16'h1);
  assign twiddle4_1_239_real = T24508 + T24506;
  assign T24506 = $signed(T24507) / $signed(22'h100000);
  assign T24507 = $signed(31'h2ad586a3) * $signed(16'h0);
  assign T24508 = $signed(T24509) / $signed(22'h100000);
  assign T24509 = $signed(31'h2f8d7139) * $signed(16'h1);
  assign T24510 = T18725[1'h0:1'h0];
  assign T24511 = T18725[1'h1:1'h1];
  assign T24512 = T18725[2'h2:2'h2];
  assign T24513 = T18725[2'h3:2'h3];
  assign T24514 = T24607 ? T24561 : T24515;
  assign T24515 = T24560 ? T24538 : T24516;
  assign T24516 = T24537 ? T24527 : T24517;
  assign T24517 = T24526 ? twiddle4_1_241_real : twiddle4_1_240_real;
  assign twiddle4_1_240_real = T24520 + T24518;
  assign T24518 = $signed(T24519) / $signed(22'h100000);
  assign T24519 = $signed(31'h2afad269) * $signed(16'h0);
  assign T24520 = $signed(T24521) / $signed(22'h100000);
  assign T24521 = $signed(31'h2f6bbe44) * $signed(16'h1);
  assign twiddle4_1_241_real = T24524 + T24522;
  assign T24522 = $signed(T24523) / $signed(22'h100000);
  assign T24523 = $signed(31'h2b2003ab) * $signed(16'h0);
  assign T24524 = $signed(T24525) / $signed(22'h100000);
  assign T24525 = $signed(31'h2f49ee0f) * $signed(16'h1);
  assign T24526 = T18725[1'h0:1'h0];
  assign T24527 = T24536 ? twiddle4_1_243_real : twiddle4_1_242_real;
  assign twiddle4_1_242_real = T24530 + T24528;
  assign T24528 = $signed(T24529) / $signed(22'h100000);
  assign T24529 = $signed(31'h2b451a54) * $signed(16'h0);
  assign T24530 = $signed(T24531) / $signed(22'h100000);
  assign T24531 = $signed(31'h2f2800ae) * $signed(16'h1);
  assign twiddle4_1_243_real = T24534 + T24532;
  assign T24532 = $signed(T24533) / $signed(22'h100000);
  assign T24533 = $signed(31'h2b6a164c) * $signed(16'h0);
  assign T24534 = $signed(T24535) / $signed(22'h100000);
  assign T24535 = $signed(31'h2f05f637) * $signed(16'h1);
  assign T24536 = T18725[1'h0:1'h0];
  assign T24537 = T18725[1'h1:1'h1];
  assign T24538 = T24559 ? T24549 : T24539;
  assign T24539 = T24548 ? twiddle4_1_245_real : twiddle4_1_244_real;
  assign twiddle4_1_244_real = T24542 + T24540;
  assign T24540 = $signed(T24541) / $signed(22'h100000);
  assign T24541 = $signed(31'h2b8ef77c) * $signed(16'h0);
  assign T24542 = $signed(T24543) / $signed(22'h100000);
  assign T24543 = $signed(31'h2ee3cebe) * $signed(16'h1);
  assign twiddle4_1_245_real = T24546 + T24544;
  assign T24544 = $signed(T24545) / $signed(22'h100000);
  assign T24545 = $signed(31'h2bb3bdce) * $signed(16'h0);
  assign T24546 = $signed(T24547) / $signed(22'h100000);
  assign T24547 = $signed(31'h2ec18a58) * $signed(16'h1);
  assign T24548 = T18725[1'h0:1'h0];
  assign T24549 = T24558 ? twiddle4_1_247_real : twiddle4_1_246_real;
  assign twiddle4_1_246_real = T24552 + T24550;
  assign T24550 = $signed(T24551) / $signed(22'h100000);
  assign T24551 = $signed(31'h2bd8692b) * $signed(16'h0);
  assign T24552 = $signed(T24553) / $signed(22'h100000);
  assign T24553 = $signed(31'h2e9f291b) * $signed(16'h1);
  assign twiddle4_1_247_real = T24556 + T24554;
  assign T24554 = $signed(T24555) / $signed(22'h100000);
  assign T24555 = $signed(31'h2bfcf97b) * $signed(16'h0);
  assign T24556 = $signed(T24557) / $signed(22'h100000);
  assign T24557 = $signed(31'h2e7cab1c) * $signed(16'h1);
  assign T24558 = T18725[1'h0:1'h0];
  assign T24559 = T18725[1'h1:1'h1];
  assign T24560 = T18725[2'h2:2'h2];
  assign T24561 = T24606 ? T24584 : T24562;
  assign T24562 = T24583 ? T24573 : T24563;
  assign T24563 = T24572 ? twiddle4_1_249_real : twiddle4_1_248_real;
  assign twiddle4_1_248_real = T24566 + T24564;
  assign T24564 = $signed(T24565) / $signed(22'h100000);
  assign T24565 = $signed(31'h2c216eaa) * $signed(16'h0);
  assign T24566 = $signed(T24567) / $signed(22'h100000);
  assign T24567 = $signed(31'h2e5a106f) * $signed(16'h1);
  assign twiddle4_1_249_real = T24570 + T24568;
  assign T24568 = $signed(T24569) / $signed(22'h100000);
  assign T24569 = $signed(31'h2c45c89f) * $signed(16'h0);
  assign T24570 = $signed(T24571) / $signed(22'h100000);
  assign T24571 = $signed(31'h2e37592c) * $signed(16'h1);
  assign T24572 = T18725[1'h0:1'h0];
  assign T24573 = T24582 ? twiddle4_1_251_real : twiddle4_1_250_real;
  assign twiddle4_1_250_real = T24576 + T24574;
  assign T24574 = $signed(T24575) / $signed(22'h100000);
  assign T24575 = $signed(31'h2c6a0746) * $signed(16'h0);
  assign T24576 = $signed(T24577) / $signed(22'h100000);
  assign T24577 = $signed(31'h2e148566) * $signed(16'h1);
  assign twiddle4_1_251_real = T24580 + T24578;
  assign T24578 = $signed(T24579) / $signed(22'h100000);
  assign T24579 = $signed(31'h2c8e2a86) * $signed(16'h0);
  assign T24580 = $signed(T24581) / $signed(22'h100000);
  assign T24581 = $signed(31'h2df19533) * $signed(16'h1);
  assign T24582 = T18725[1'h0:1'h0];
  assign T24583 = T18725[1'h1:1'h1];
  assign T24584 = T24605 ? T24595 : T24585;
  assign T24585 = T24594 ? twiddle4_1_253_real : twiddle4_1_252_real;
  assign twiddle4_1_252_real = T24588 + T24586;
  assign T24586 = $signed(T24587) / $signed(22'h100000);
  assign T24587 = $signed(31'h2cb2324b) * $signed(16'h0);
  assign T24588 = $signed(T24589) / $signed(22'h100000);
  assign T24589 = $signed(31'h2dce88a9) * $signed(16'h1);
  assign twiddle4_1_253_real = T24592 + T24590;
  assign T24590 = $signed(T24591) / $signed(22'h100000);
  assign T24591 = $signed(31'h2cd61e7e) * $signed(16'h0);
  assign T24592 = $signed(T24593) / $signed(22'h100000);
  assign T24593 = $signed(31'h2dab5fde) * $signed(16'h1);
  assign T24594 = T18725[1'h0:1'h0];
  assign T24595 = T24604 ? twiddle4_1_255_real : twiddle4_1_254_real;
  assign twiddle4_1_254_real = T24598 + T24596;
  assign T24596 = $signed(T24597) / $signed(22'h100000);
  assign T24597 = $signed(31'h2cf9ef09) * $signed(16'h0);
  assign T24598 = $signed(T24599) / $signed(22'h100000);
  assign T24599 = $signed(31'h2d881ae7) * $signed(16'h1);
  assign twiddle4_1_255_real = T24602 + T24600;
  assign T24600 = $signed(T24601) / $signed(22'h100000);
  assign T24601 = $signed(31'h2d1da3d5) * $signed(16'h0);
  assign T24602 = $signed(T24603) / $signed(22'h100000);
  assign T24603 = $signed(31'h2d64b9da) * $signed(16'h1);
  assign T24604 = T18725[1'h0:1'h0];
  assign T24605 = T18725[1'h1:1'h1];
  assign T24606 = T18725[2'h2:2'h2];
  assign T24607 = T18725[2'h3:2'h3];
  assign T24608 = T18725[3'h4:3'h4];
  assign T24609 = T18725[3'h5:3'h5];
  assign T24610 = T18725[3'h6:3'h6];
  assign T24611 = T23759[6'h2e:6'h2e];
  assign T24612 = T18725[3'h7:3'h7];
  assign T24613 = {T26570, T24614};
  assign T24614 = T26569 ? T25465 : T24615;
  assign T24615 = T25464 ? T24998 : T24616;
  assign T24616 = T24997 ? T24807 : T24617;
  assign T24617 = T24806 ? T24712 : T24618;
  assign T24618 = T24711 ? T24665 : T24619;
  assign T24619 = T24664 ? T24642 : T24620;
  assign T24620 = T24641 ? T24631 : T24621;
  assign T24621 = T24630 ? twiddle4_1_257_real : twiddle4_1_256_real;
  assign twiddle4_1_256_real = T24624 + T24622;
  assign T24622 = $signed(T24623) / $signed(22'h100000);
  assign T24623 = $signed(31'h2d413ccc) * $signed(16'h0);
  assign T24624 = $signed(T24625) / $signed(22'h100000);
  assign T24625 = $signed(31'h2d413ccc) * $signed(16'h1);
  assign twiddle4_1_257_real = T24628 + T24626;
  assign T24626 = $signed(T24627) / $signed(22'h100000);
  assign T24627 = $signed(31'h2d64b9da) * $signed(16'h0);
  assign T24628 = $signed(T24629) / $signed(22'h100000);
  assign T24629 = $signed(31'h2d1da3d5) * $signed(16'h1);
  assign T24630 = T18725[1'h0:1'h0];
  assign T24631 = T24640 ? twiddle4_1_259_real : twiddle4_1_258_real;
  assign twiddle4_1_258_real = T24634 + T24632;
  assign T24632 = $signed(T24633) / $signed(22'h100000);
  assign T24633 = $signed(31'h2d881ae7) * $signed(16'h0);
  assign T24634 = $signed(T24635) / $signed(22'h100000);
  assign T24635 = $signed(31'h2cf9ef09) * $signed(16'h1);
  assign twiddle4_1_259_real = T24638 + T24636;
  assign T24636 = $signed(T24637) / $signed(22'h100000);
  assign T24637 = $signed(31'h2dab5fde) * $signed(16'h0);
  assign T24638 = $signed(T24639) / $signed(22'h100000);
  assign T24639 = $signed(31'h2cd61e7e) * $signed(16'h1);
  assign T24640 = T18725[1'h0:1'h0];
  assign T24641 = T18725[1'h1:1'h1];
  assign T24642 = T24663 ? T24653 : T24643;
  assign T24643 = T24652 ? twiddle4_1_261_real : twiddle4_1_260_real;
  assign twiddle4_1_260_real = T24646 + T24644;
  assign T24644 = $signed(T24645) / $signed(22'h100000);
  assign T24645 = $signed(31'h2dce88a9) * $signed(16'h0);
  assign T24646 = $signed(T24647) / $signed(22'h100000);
  assign T24647 = $signed(31'h2cb2324b) * $signed(16'h1);
  assign twiddle4_1_261_real = T24650 + T24648;
  assign T24648 = $signed(T24649) / $signed(22'h100000);
  assign T24649 = $signed(31'h2df19533) * $signed(16'h0);
  assign T24650 = $signed(T24651) / $signed(22'h100000);
  assign T24651 = $signed(31'h2c8e2a86) * $signed(16'h1);
  assign T24652 = T18725[1'h0:1'h0];
  assign T24653 = T24662 ? twiddle4_1_263_real : twiddle4_1_262_real;
  assign twiddle4_1_262_real = T24656 + T24654;
  assign T24654 = $signed(T24655) / $signed(22'h100000);
  assign T24655 = $signed(31'h2e148566) * $signed(16'h0);
  assign T24656 = $signed(T24657) / $signed(22'h100000);
  assign T24657 = $signed(31'h2c6a0746) * $signed(16'h1);
  assign twiddle4_1_263_real = T24660 + T24658;
  assign T24658 = $signed(T24659) / $signed(22'h100000);
  assign T24659 = $signed(31'h2e37592c) * $signed(16'h0);
  assign T24660 = $signed(T24661) / $signed(22'h100000);
  assign T24661 = $signed(31'h2c45c89f) * $signed(16'h1);
  assign T24662 = T18725[1'h0:1'h0];
  assign T24663 = T18725[1'h1:1'h1];
  assign T24664 = T18725[2'h2:2'h2];
  assign T24665 = T24710 ? T24688 : T24666;
  assign T24666 = T24687 ? T24677 : T24667;
  assign T24667 = T24676 ? twiddle4_1_265_real : twiddle4_1_264_real;
  assign twiddle4_1_264_real = T24670 + T24668;
  assign T24668 = $signed(T24669) / $signed(22'h100000);
  assign T24669 = $signed(31'h2e5a106f) * $signed(16'h0);
  assign T24670 = $signed(T24671) / $signed(22'h100000);
  assign T24671 = $signed(31'h2c216eaa) * $signed(16'h1);
  assign twiddle4_1_265_real = T24674 + T24672;
  assign T24672 = $signed(T24673) / $signed(22'h100000);
  assign T24673 = $signed(31'h2e7cab1c) * $signed(16'h0);
  assign T24674 = $signed(T24675) / $signed(22'h100000);
  assign T24675 = $signed(31'h2bfcf97b) * $signed(16'h1);
  assign T24676 = T18725[1'h0:1'h0];
  assign T24677 = T24686 ? twiddle4_1_267_real : twiddle4_1_266_real;
  assign twiddle4_1_266_real = T24680 + T24678;
  assign T24678 = $signed(T24679) / $signed(22'h100000);
  assign T24679 = $signed(31'h2e9f291b) * $signed(16'h0);
  assign T24680 = $signed(T24681) / $signed(22'h100000);
  assign T24681 = $signed(31'h2bd8692b) * $signed(16'h1);
  assign twiddle4_1_267_real = T24684 + T24682;
  assign T24682 = $signed(T24683) / $signed(22'h100000);
  assign T24683 = $signed(31'h2ec18a58) * $signed(16'h0);
  assign T24684 = $signed(T24685) / $signed(22'h100000);
  assign T24685 = $signed(31'h2bb3bdce) * $signed(16'h1);
  assign T24686 = T18725[1'h0:1'h0];
  assign T24687 = T18725[1'h1:1'h1];
  assign T24688 = T24709 ? T24699 : T24689;
  assign T24689 = T24698 ? twiddle4_1_269_real : twiddle4_1_268_real;
  assign twiddle4_1_268_real = T24692 + T24690;
  assign T24690 = $signed(T24691) / $signed(22'h100000);
  assign T24691 = $signed(31'h2ee3cebe) * $signed(16'h0);
  assign T24692 = $signed(T24693) / $signed(22'h100000);
  assign T24693 = $signed(31'h2b8ef77c) * $signed(16'h1);
  assign twiddle4_1_269_real = T24696 + T24694;
  assign T24694 = $signed(T24695) / $signed(22'h100000);
  assign T24695 = $signed(31'h2f05f637) * $signed(16'h0);
  assign T24696 = $signed(T24697) / $signed(22'h100000);
  assign T24697 = $signed(31'h2b6a164c) * $signed(16'h1);
  assign T24698 = T18725[1'h0:1'h0];
  assign T24699 = T24708 ? twiddle4_1_271_real : twiddle4_1_270_real;
  assign twiddle4_1_270_real = T24702 + T24700;
  assign T24700 = $signed(T24701) / $signed(22'h100000);
  assign T24701 = $signed(31'h2f2800ae) * $signed(16'h0);
  assign T24702 = $signed(T24703) / $signed(22'h100000);
  assign T24703 = $signed(31'h2b451a54) * $signed(16'h1);
  assign twiddle4_1_271_real = T24706 + T24704;
  assign T24704 = $signed(T24705) / $signed(22'h100000);
  assign T24705 = $signed(31'h2f49ee0f) * $signed(16'h0);
  assign T24706 = $signed(T24707) / $signed(22'h100000);
  assign T24707 = $signed(31'h2b2003ab) * $signed(16'h1);
  assign T24708 = T18725[1'h0:1'h0];
  assign T24709 = T18725[1'h1:1'h1];
  assign T24710 = T18725[2'h2:2'h2];
  assign T24711 = T18725[2'h3:2'h3];
  assign T24712 = T24805 ? T24759 : T24713;
  assign T24713 = T24758 ? T24736 : T24714;
  assign T24714 = T24735 ? T24725 : T24715;
  assign T24715 = T24724 ? twiddle4_1_273_real : twiddle4_1_272_real;
  assign twiddle4_1_272_real = T24718 + T24716;
  assign T24716 = $signed(T24717) / $signed(22'h100000);
  assign T24717 = $signed(31'h2f6bbe44) * $signed(16'h0);
  assign T24718 = $signed(T24719) / $signed(22'h100000);
  assign T24719 = $signed(31'h2afad269) * $signed(16'h1);
  assign twiddle4_1_273_real = T24722 + T24720;
  assign T24720 = $signed(T24721) / $signed(22'h100000);
  assign T24721 = $signed(31'h2f8d7139) * $signed(16'h0);
  assign T24722 = $signed(T24723) / $signed(22'h100000);
  assign T24723 = $signed(31'h2ad586a3) * $signed(16'h1);
  assign T24724 = T18725[1'h0:1'h0];
  assign T24725 = T24734 ? twiddle4_1_275_real : twiddle4_1_274_real;
  assign twiddle4_1_274_real = T24728 + T24726;
  assign T24726 = $signed(T24727) / $signed(22'h100000);
  assign T24727 = $signed(31'h2faf06d9) * $signed(16'h0);
  assign T24728 = $signed(T24729) / $signed(22'h100000);
  assign T24729 = $signed(31'h2ab02071) * $signed(16'h1);
  assign twiddle4_1_275_real = T24732 + T24730;
  assign T24730 = $signed(T24731) / $signed(22'h100000);
  assign T24731 = $signed(31'h2fd07f0f) * $signed(16'h0);
  assign T24732 = $signed(T24733) / $signed(22'h100000);
  assign T24733 = $signed(31'h2a8a9fea) * $signed(16'h1);
  assign T24734 = T18725[1'h0:1'h0];
  assign T24735 = T18725[1'h1:1'h1];
  assign T24736 = T24757 ? T24747 : T24737;
  assign T24737 = T24746 ? twiddle4_1_277_real : twiddle4_1_276_real;
  assign twiddle4_1_276_real = T24740 + T24738;
  assign T24738 = $signed(T24739) / $signed(22'h100000);
  assign T24739 = $signed(31'h2ff1d9c6) * $signed(16'h0);
  assign T24740 = $signed(T24741) / $signed(22'h100000);
  assign T24741 = $signed(31'h2a650525) * $signed(16'h1);
  assign twiddle4_1_277_real = T24744 + T24742;
  assign T24742 = $signed(T24743) / $signed(22'h100000);
  assign T24743 = $signed(31'h301316ea) * $signed(16'h0);
  assign T24744 = $signed(T24745) / $signed(22'h100000);
  assign T24745 = $signed(31'h2a3f5039) * $signed(16'h1);
  assign T24746 = T18725[1'h0:1'h0];
  assign T24747 = T24756 ? twiddle4_1_279_real : twiddle4_1_278_real;
  assign twiddle4_1_278_real = T24750 + T24748;
  assign T24748 = $signed(T24749) / $signed(22'h100000);
  assign T24749 = $signed(31'h30343667) * $signed(16'h0);
  assign T24750 = $signed(T24751) / $signed(22'h100000);
  assign T24751 = $signed(31'h2a19813e) * $signed(16'h1);
  assign twiddle4_1_279_real = T24754 + T24752;
  assign T24752 = $signed(T24753) / $signed(22'h100000);
  assign T24753 = $signed(31'h30553827) * $signed(16'h0);
  assign T24754 = $signed(T24755) / $signed(22'h100000);
  assign T24755 = $signed(31'h29f3984b) * $signed(16'h1);
  assign T24756 = T18725[1'h0:1'h0];
  assign T24757 = T18725[1'h1:1'h1];
  assign T24758 = T18725[2'h2:2'h2];
  assign T24759 = T24804 ? T24782 : T24760;
  assign T24760 = T24781 ? T24771 : T24761;
  assign T24761 = T24770 ? twiddle4_1_281_real : twiddle4_1_280_real;
  assign twiddle4_1_280_real = T24764 + T24762;
  assign T24762 = $signed(T24763) / $signed(22'h100000);
  assign T24763 = $signed(31'h30761c17) * $signed(16'h0);
  assign T24764 = $signed(T24765) / $signed(22'h100000);
  assign T24765 = $signed(31'h29cd9577) * $signed(16'h1);
  assign twiddle4_1_281_real = T24768 + T24766;
  assign T24766 = $signed(T24767) / $signed(22'h100000);
  assign T24767 = $signed(31'h3096e223) * $signed(16'h0);
  assign T24768 = $signed(T24769) / $signed(22'h100000);
  assign T24769 = $signed(31'h29a778da) * $signed(16'h1);
  assign T24770 = T18725[1'h0:1'h0];
  assign T24771 = T24780 ? twiddle4_1_283_real : twiddle4_1_282_real;
  assign twiddle4_1_282_real = T24774 + T24772;
  assign T24772 = $signed(T24773) / $signed(22'h100000);
  assign T24773 = $signed(31'h30b78a35) * $signed(16'h0);
  assign T24774 = $signed(T24775) / $signed(22'h100000);
  assign T24775 = $signed(31'h2981428b) * $signed(16'h1);
  assign twiddle4_1_283_real = T24778 + T24776;
  assign T24776 = $signed(T24777) / $signed(22'h100000);
  assign T24777 = $signed(31'h30d8143b) * $signed(16'h0);
  assign T24778 = $signed(T24779) / $signed(22'h100000);
  assign T24779 = $signed(31'h295af2a2) * $signed(16'h1);
  assign T24780 = T18725[1'h0:1'h0];
  assign T24781 = T18725[1'h1:1'h1];
  assign T24782 = T24803 ? T24793 : T24783;
  assign T24783 = T24792 ? twiddle4_1_285_real : twiddle4_1_284_real;
  assign twiddle4_1_284_real = T24786 + T24784;
  assign T24784 = $signed(T24785) / $signed(22'h100000);
  assign T24785 = $signed(31'h30f8801f) * $signed(16'h0);
  assign T24786 = $signed(T24787) / $signed(22'h100000);
  assign T24787 = $signed(31'h29348937) * $signed(16'h1);
  assign twiddle4_1_285_real = T24790 + T24788;
  assign T24788 = $signed(T24789) / $signed(22'h100000);
  assign T24789 = $signed(31'h3118cdce) * $signed(16'h0);
  assign T24790 = $signed(T24791) / $signed(22'h100000);
  assign T24791 = $signed(31'h290e0660) * $signed(16'h1);
  assign T24792 = T18725[1'h0:1'h0];
  assign T24793 = T24802 ? twiddle4_1_287_real : twiddle4_1_286_real;
  assign twiddle4_1_286_real = T24796 + T24794;
  assign T24794 = $signed(T24795) / $signed(22'h100000);
  assign T24795 = $signed(31'h3138fd34) * $signed(16'h0);
  assign T24796 = $signed(T24797) / $signed(22'h100000);
  assign T24797 = $signed(31'h28e76a37) * $signed(16'h1);
  assign twiddle4_1_287_real = T24800 + T24798;
  assign T24798 = $signed(T24799) / $signed(22'h100000);
  assign T24799 = $signed(31'h31590e3d) * $signed(16'h0);
  assign T24800 = $signed(T24801) / $signed(22'h100000);
  assign T24801 = $signed(31'h28c0b4d2) * $signed(16'h1);
  assign T24802 = T18725[1'h0:1'h0];
  assign T24803 = T18725[1'h1:1'h1];
  assign T24804 = T18725[2'h2:2'h2];
  assign T24805 = T18725[2'h3:2'h3];
  assign T24806 = T18725[3'h4:3'h4];
  assign T24807 = T24996 ? T24902 : T24808;
  assign T24808 = T24901 ? T24855 : T24809;
  assign T24809 = T24854 ? T24832 : T24810;
  assign T24810 = T24831 ? T24821 : T24811;
  assign T24811 = T24820 ? twiddle4_1_289_real : twiddle4_1_288_real;
  assign twiddle4_1_288_real = T24814 + T24812;
  assign T24812 = $signed(T24813) / $signed(22'h100000);
  assign T24813 = $signed(31'h317900d6) * $signed(16'h0);
  assign T24814 = $signed(T24815) / $signed(22'h100000);
  assign T24815 = $signed(31'h2899e64a) * $signed(16'h1);
  assign twiddle4_1_289_real = T24818 + T24816;
  assign T24816 = $signed(T24817) / $signed(22'h100000);
  assign T24817 = $signed(31'h3198d4ea) * $signed(16'h0);
  assign T24818 = $signed(T24819) / $signed(22'h100000);
  assign T24819 = $signed(31'h2872feb6) * $signed(16'h1);
  assign T24820 = T18725[1'h0:1'h0];
  assign T24821 = T24830 ? twiddle4_1_291_real : twiddle4_1_290_real;
  assign twiddle4_1_290_real = T24824 + T24822;
  assign T24822 = $signed(T24823) / $signed(22'h100000);
  assign T24823 = $signed(31'h31b88a66) * $signed(16'h0);
  assign T24824 = $signed(T24825) / $signed(22'h100000);
  assign T24825 = $signed(31'h284bfe2f) * $signed(16'h1);
  assign twiddle4_1_291_real = T24828 + T24826;
  assign T24826 = $signed(T24827) / $signed(22'h100000);
  assign T24827 = $signed(31'h31d82136) * $signed(16'h0);
  assign T24828 = $signed(T24829) / $signed(22'h100000);
  assign T24829 = $signed(31'h2824e4cc) * $signed(16'h1);
  assign T24830 = T18725[1'h0:1'h0];
  assign T24831 = T18725[1'h1:1'h1];
  assign T24832 = T24853 ? T24843 : T24833;
  assign T24833 = T24842 ? twiddle4_1_293_real : twiddle4_1_292_real;
  assign twiddle4_1_292_real = T24836 + T24834;
  assign T24834 = $signed(T24835) / $signed(22'h100000);
  assign T24835 = $signed(31'h31f79947) * $signed(16'h0);
  assign T24836 = $signed(T24837) / $signed(22'h100000);
  assign T24837 = $signed(31'h27fdb2a6) * $signed(16'h1);
  assign twiddle4_1_293_real = T24840 + T24838;
  assign T24838 = $signed(T24839) / $signed(22'h100000);
  assign T24839 = $signed(31'h3216f286) * $signed(16'h0);
  assign T24840 = $signed(T24841) / $signed(22'h100000);
  assign T24841 = $signed(31'h27d667d5) * $signed(16'h1);
  assign T24842 = T18725[1'h0:1'h0];
  assign T24843 = T24852 ? twiddle4_1_295_real : twiddle4_1_294_real;
  assign twiddle4_1_294_real = T24846 + T24844;
  assign T24844 = $signed(T24845) / $signed(22'h100000);
  assign T24845 = $signed(31'h32362cdf) * $signed(16'h0);
  assign T24846 = $signed(T24847) / $signed(22'h100000);
  assign T24847 = $signed(31'h27af0471) * $signed(16'h1);
  assign twiddle4_1_295_real = T24850 + T24848;
  assign T24848 = $signed(T24849) / $signed(22'h100000);
  assign T24849 = $signed(31'h3255483f) * $signed(16'h0);
  assign T24850 = $signed(T24851) / $signed(22'h100000);
  assign T24851 = $signed(31'h27878893) * $signed(16'h1);
  assign T24852 = T18725[1'h0:1'h0];
  assign T24853 = T18725[1'h1:1'h1];
  assign T24854 = T18725[2'h2:2'h2];
  assign T24855 = T24900 ? T24878 : T24856;
  assign T24856 = T24877 ? T24867 : T24857;
  assign T24857 = T24866 ? twiddle4_1_297_real : twiddle4_1_296_real;
  assign twiddle4_1_296_real = T24860 + T24858;
  assign T24858 = $signed(T24859) / $signed(22'h100000);
  assign T24859 = $signed(31'h32744493) * $signed(16'h0);
  assign T24860 = $signed(T24861) / $signed(22'h100000);
  assign T24861 = $signed(31'h275ff452) * $signed(16'h1);
  assign twiddle4_1_297_real = T24864 + T24862;
  assign T24862 = $signed(T24863) / $signed(22'h100000);
  assign T24863 = $signed(31'h329321c7) * $signed(16'h0);
  assign T24864 = $signed(T24865) / $signed(22'h100000);
  assign T24865 = $signed(31'h273847c7) * $signed(16'h1);
  assign T24866 = T18725[1'h0:1'h0];
  assign T24867 = T24876 ? twiddle4_1_299_real : twiddle4_1_298_real;
  assign twiddle4_1_298_real = T24870 + T24868;
  assign T24868 = $signed(T24869) / $signed(22'h100000);
  assign T24869 = $signed(31'h32b1dfc9) * $signed(16'h0);
  assign T24870 = $signed(T24871) / $signed(22'h100000);
  assign T24871 = $signed(31'h2710830b) * $signed(16'h1);
  assign twiddle4_1_299_real = T24874 + T24872;
  assign T24872 = $signed(T24873) / $signed(22'h100000);
  assign T24873 = $signed(31'h32d07e85) * $signed(16'h0);
  assign T24874 = $signed(T24875) / $signed(22'h100000);
  assign T24875 = $signed(31'h26e8a637) * $signed(16'h1);
  assign T24876 = T18725[1'h0:1'h0];
  assign T24877 = T18725[1'h1:1'h1];
  assign T24878 = T24899 ? T24889 : T24879;
  assign T24879 = T24888 ? twiddle4_1_301_real : twiddle4_1_300_real;
  assign twiddle4_1_300_real = T24882 + T24880;
  assign T24880 = $signed(T24881) / $signed(22'h100000);
  assign T24881 = $signed(31'h32eefde9) * $signed(16'h0);
  assign T24882 = $signed(T24883) / $signed(22'h100000);
  assign T24883 = $signed(31'h26c0b162) * $signed(16'h1);
  assign twiddle4_1_301_real = T24886 + T24884;
  assign T24884 = $signed(T24885) / $signed(22'h100000);
  assign T24885 = $signed(31'h330d5de2) * $signed(16'h0);
  assign T24886 = $signed(T24887) / $signed(22'h100000);
  assign T24887 = $signed(31'h2698a4a5) * $signed(16'h1);
  assign T24888 = T18725[1'h0:1'h0];
  assign T24889 = T24898 ? twiddle4_1_303_real : twiddle4_1_302_real;
  assign twiddle4_1_302_real = T24892 + T24890;
  assign T24890 = $signed(T24891) / $signed(22'h100000);
  assign T24891 = $signed(31'h332b9e5d) * $signed(16'h0);
  assign T24892 = $signed(T24893) / $signed(22'h100000);
  assign T24893 = $signed(31'h2670801a) * $signed(16'h1);
  assign twiddle4_1_303_real = T24896 + T24894;
  assign T24894 = $signed(T24895) / $signed(22'h100000);
  assign T24895 = $signed(31'h3349bf48) * $signed(16'h0);
  assign T24896 = $signed(T24897) / $signed(22'h100000);
  assign T24897 = $signed(31'h264843d8) * $signed(16'h1);
  assign T24898 = T18725[1'h0:1'h0];
  assign T24899 = T18725[1'h1:1'h1];
  assign T24900 = T18725[2'h2:2'h2];
  assign T24901 = T18725[2'h3:2'h3];
  assign T24902 = T24995 ? T24949 : T24903;
  assign T24903 = T24948 ? T24926 : T24904;
  assign T24904 = T24925 ? T24915 : T24905;
  assign T24905 = T24914 ? twiddle4_1_305_real : twiddle4_1_304_real;
  assign twiddle4_1_304_real = T24908 + T24906;
  assign T24906 = $signed(T24907) / $signed(22'h100000);
  assign T24907 = $signed(31'h3367c08f) * $signed(16'h0);
  assign T24908 = $signed(T24909) / $signed(22'h100000);
  assign T24909 = $signed(31'h261feff9) * $signed(16'h1);
  assign twiddle4_1_305_real = T24912 + T24910;
  assign T24910 = $signed(T24911) / $signed(22'h100000);
  assign T24911 = $signed(31'h3385a221) * $signed(16'h0);
  assign T24912 = $signed(T24913) / $signed(22'h100000);
  assign T24913 = $signed(31'h25f78496) * $signed(16'h1);
  assign T24914 = T18725[1'h0:1'h0];
  assign T24915 = T24924 ? twiddle4_1_307_real : twiddle4_1_306_real;
  assign twiddle4_1_306_real = T24918 + T24916;
  assign T24916 = $signed(T24917) / $signed(22'h100000);
  assign T24917 = $signed(31'h33a363eb) * $signed(16'h0);
  assign T24918 = $signed(T24919) / $signed(22'h100000);
  assign T24919 = $signed(31'h25cf01c7) * $signed(16'h1);
  assign twiddle4_1_307_real = T24922 + T24920;
  assign T24920 = $signed(T24921) / $signed(22'h100000);
  assign T24921 = $signed(31'h33c105db) * $signed(16'h0);
  assign T24922 = $signed(T24923) / $signed(22'h100000);
  assign T24923 = $signed(31'h25a667a6) * $signed(16'h1);
  assign T24924 = T18725[1'h0:1'h0];
  assign T24925 = T18725[1'h1:1'h1];
  assign T24926 = T24947 ? T24937 : T24927;
  assign T24927 = T24936 ? twiddle4_1_309_real : twiddle4_1_308_real;
  assign twiddle4_1_308_real = T24930 + T24928;
  assign T24928 = $signed(T24929) / $signed(22'h100000);
  assign T24929 = $signed(31'h33de87de) * $signed(16'h0);
  assign T24930 = $signed(T24931) / $signed(22'h100000);
  assign T24931 = $signed(31'h257db64b) * $signed(16'h1);
  assign twiddle4_1_309_real = T24934 + T24932;
  assign T24932 = $signed(T24933) / $signed(22'h100000);
  assign T24933 = $signed(31'h33fbe9e2) * $signed(16'h0);
  assign T24934 = $signed(T24935) / $signed(22'h100000);
  assign T24935 = $signed(31'h2554edd0) * $signed(16'h1);
  assign T24936 = T18725[1'h0:1'h0];
  assign T24937 = T24946 ? twiddle4_1_311_real : twiddle4_1_310_real;
  assign twiddle4_1_310_real = T24940 + T24938;
  assign T24938 = $signed(T24939) / $signed(22'h100000);
  assign T24939 = $signed(31'h34192bd5) * $signed(16'h0);
  assign T24940 = $signed(T24941) / $signed(22'h100000);
  assign T24941 = $signed(31'h252c0e4e) * $signed(16'h1);
  assign twiddle4_1_311_real = T24944 + T24942;
  assign T24942 = $signed(T24943) / $signed(22'h100000);
  assign T24943 = $signed(31'h34364da5) * $signed(16'h0);
  assign T24944 = $signed(T24945) / $signed(22'h100000);
  assign T24945 = $signed(31'h250317de) * $signed(16'h1);
  assign T24946 = T18725[1'h0:1'h0];
  assign T24947 = T18725[1'h1:1'h1];
  assign T24948 = T18725[2'h2:2'h2];
  assign T24949 = T24994 ? T24972 : T24950;
  assign T24950 = T24971 ? T24961 : T24951;
  assign T24951 = T24960 ? twiddle4_1_313_real : twiddle4_1_312_real;
  assign twiddle4_1_312_real = T24954 + T24952;
  assign T24952 = $signed(T24953) / $signed(22'h100000);
  assign T24953 = $signed(31'h34534f40) * $signed(16'h0);
  assign T24954 = $signed(T24955) / $signed(22'h100000);
  assign T24955 = $signed(31'h24da0a99) * $signed(16'h1);
  assign twiddle4_1_313_real = T24958 + T24956;
  assign T24956 = $signed(T24957) / $signed(22'h100000);
  assign T24957 = $signed(31'h34703094) * $signed(16'h0);
  assign T24958 = $signed(T24959) / $signed(22'h100000);
  assign T24959 = $signed(31'h24b0e699) * $signed(16'h1);
  assign T24960 = T18725[1'h0:1'h0];
  assign T24961 = T24970 ? twiddle4_1_315_real : twiddle4_1_314_real;
  assign twiddle4_1_314_real = T24964 + T24962;
  assign T24962 = $signed(T24963) / $signed(22'h100000);
  assign T24963 = $signed(31'h348cf190) * $signed(16'h0);
  assign T24964 = $signed(T24965) / $signed(22'h100000);
  assign T24965 = $signed(31'h2487abf7) * $signed(16'h1);
  assign twiddle4_1_315_real = T24968 + T24966;
  assign T24966 = $signed(T24967) / $signed(22'h100000);
  assign T24967 = $signed(31'h34a99221) * $signed(16'h0);
  assign T24968 = $signed(T24969) / $signed(22'h100000);
  assign T24969 = $signed(31'h245e5acc) * $signed(16'h1);
  assign T24970 = T18725[1'h0:1'h0];
  assign T24971 = T18725[1'h1:1'h1];
  assign T24972 = T24993 ? T24983 : T24973;
  assign T24973 = T24982 ? twiddle4_1_317_real : twiddle4_1_316_real;
  assign twiddle4_1_316_real = T24976 + T24974;
  assign T24974 = $signed(T24975) / $signed(22'h100000);
  assign T24975 = $signed(31'h34c61236) * $signed(16'h0);
  assign T24976 = $signed(T24977) / $signed(22'h100000);
  assign T24977 = $signed(31'h2434f332) * $signed(16'h1);
  assign twiddle4_1_317_real = T24980 + T24978;
  assign T24978 = $signed(T24979) / $signed(22'h100000);
  assign T24979 = $signed(31'h34e271bd) * $signed(16'h0);
  assign T24980 = $signed(T24981) / $signed(22'h100000);
  assign T24981 = $signed(31'h240b7542) * $signed(16'h1);
  assign T24982 = T18725[1'h0:1'h0];
  assign T24983 = T24992 ? twiddle4_1_319_real : twiddle4_1_318_real;
  assign twiddle4_1_318_real = T24986 + T24984;
  assign T24984 = $signed(T24985) / $signed(22'h100000);
  assign T24985 = $signed(31'h34feb0a5) * $signed(16'h0);
  assign T24986 = $signed(T24987) / $signed(22'h100000);
  assign T24987 = $signed(31'h23e1e117) * $signed(16'h1);
  assign twiddle4_1_319_real = T24990 + T24988;
  assign T24988 = $signed(T24989) / $signed(22'h100000);
  assign T24989 = $signed(31'h351acedc) * $signed(16'h0);
  assign T24990 = $signed(T24991) / $signed(22'h100000);
  assign T24991 = $signed(31'h23b836c9) * $signed(16'h1);
  assign T24992 = T18725[1'h0:1'h0];
  assign T24993 = T18725[1'h1:1'h1];
  assign T24994 = T18725[2'h2:2'h2];
  assign T24995 = T18725[2'h3:2'h3];
  assign T24996 = T18725[3'h4:3'h4];
  assign T24997 = T18725[3'h5:3'h5];
  assign T24998 = T25463 ? T25209 : T24999;
  assign T24999 = T25208 ? T25094 : T25000;
  assign T25000 = T25093 ? T25047 : T25001;
  assign T25001 = T25046 ? T25024 : T25002;
  assign T25002 = T25023 ? T25013 : T25003;
  assign T25003 = T25012 ? twiddle4_1_321_real : twiddle4_1_320_real;
  assign twiddle4_1_320_real = T25006 + T25004;
  assign T25004 = $signed(T25005) / $signed(22'h100000);
  assign T25005 = $signed(31'h3536cc52) * $signed(16'h0);
  assign T25006 = $signed(T25007) / $signed(22'h100000);
  assign T25007 = $signed(31'h238e7673) * $signed(16'h1);
  assign twiddle4_1_321_real = T25010 + T25008;
  assign T25008 = $signed(T25009) / $signed(22'h100000);
  assign T25009 = $signed(31'h3552a8f4) * $signed(16'h0);
  assign T25010 = $signed(T25011) / $signed(22'h100000);
  assign T25011 = $signed(31'h2364a02e) * $signed(16'h1);
  assign T25012 = T18725[1'h0:1'h0];
  assign T25013 = T25022 ? twiddle4_1_323_real : twiddle4_1_322_real;
  assign twiddle4_1_322_real = T25016 + T25014;
  assign T25014 = $signed(T25015) / $signed(22'h100000);
  assign T25015 = $signed(31'h356e64b2) * $signed(16'h0);
  assign T25016 = $signed(T25017) / $signed(22'h100000);
  assign T25017 = $signed(31'h233ab413) * $signed(16'h1);
  assign twiddle4_1_323_real = T25020 + T25018;
  assign T25018 = $signed(T25019) / $signed(22'h100000);
  assign T25019 = $signed(31'h3589ff7a) * $signed(16'h0);
  assign T25020 = $signed(T25021) / $signed(22'h100000);
  assign T25021 = $signed(31'h2310b23e) * $signed(16'h1);
  assign T25022 = T18725[1'h0:1'h0];
  assign T25023 = T18725[1'h1:1'h1];
  assign T25024 = T25045 ? T25035 : T25025;
  assign T25025 = T25034 ? twiddle4_1_325_real : twiddle4_1_324_real;
  assign twiddle4_1_324_real = T25028 + T25026;
  assign T25026 = $signed(T25027) / $signed(22'h100000);
  assign T25027 = $signed(31'h35a5793c) * $signed(16'h0);
  assign T25028 = $signed(T25029) / $signed(22'h100000);
  assign T25029 = $signed(31'h22e69ac7) * $signed(16'h1);
  assign twiddle4_1_325_real = T25032 + T25030;
  assign T25030 = $signed(T25031) / $signed(22'h100000);
  assign T25031 = $signed(31'h35c0d1e6) * $signed(16'h0);
  assign T25032 = $signed(T25033) / $signed(22'h100000);
  assign T25033 = $signed(31'h22bc6dc9) * $signed(16'h1);
  assign T25034 = T18725[1'h0:1'h0];
  assign T25035 = T25044 ? twiddle4_1_327_real : twiddle4_1_326_real;
  assign twiddle4_1_326_real = T25038 + T25036;
  assign T25036 = $signed(T25037) / $signed(22'h100000);
  assign T25037 = $signed(31'h35dc0968) * $signed(16'h0);
  assign T25038 = $signed(T25039) / $signed(22'h100000);
  assign T25039 = $signed(31'h22922b5e) * $signed(16'h1);
  assign twiddle4_1_327_real = T25042 + T25040;
  assign T25040 = $signed(T25041) / $signed(22'h100000);
  assign T25041 = $signed(31'h35f71fb1) * $signed(16'h0);
  assign T25042 = $signed(T25043) / $signed(22'h100000);
  assign T25043 = $signed(31'h2267d39f) * $signed(16'h1);
  assign T25044 = T18725[1'h0:1'h0];
  assign T25045 = T18725[1'h1:1'h1];
  assign T25046 = T18725[2'h2:2'h2];
  assign T25047 = T25092 ? T25070 : T25048;
  assign T25048 = T25069 ? T25059 : T25049;
  assign T25049 = T25058 ? twiddle4_1_329_real : twiddle4_1_328_real;
  assign twiddle4_1_328_real = T25052 + T25050;
  assign T25050 = $signed(T25051) / $signed(22'h100000);
  assign T25051 = $signed(31'h361214b0) * $signed(16'h0);
  assign T25052 = $signed(T25053) / $signed(22'h100000);
  assign T25053 = $signed(31'h223d66a8) * $signed(16'h1);
  assign twiddle4_1_329_real = T25056 + T25054;
  assign T25054 = $signed(T25055) / $signed(22'h100000);
  assign T25055 = $signed(31'h362ce854) * $signed(16'h0);
  assign T25056 = $signed(T25057) / $signed(22'h100000);
  assign T25057 = $signed(31'h2212e491) * $signed(16'h1);
  assign T25058 = T18725[1'h0:1'h0];
  assign T25059 = T25068 ? twiddle4_1_331_real : twiddle4_1_330_real;
  assign twiddle4_1_330_real = T25062 + T25060;
  assign T25060 = $signed(T25061) / $signed(22'h100000);
  assign T25061 = $signed(31'h36479a8e) * $signed(16'h0);
  assign T25062 = $signed(T25063) / $signed(22'h100000);
  assign T25063 = $signed(31'h21e84d76) * $signed(16'h1);
  assign twiddle4_1_331_real = T25066 + T25064;
  assign T25064 = $signed(T25065) / $signed(22'h100000);
  assign T25065 = $signed(31'h36622b4b) * $signed(16'h0);
  assign T25066 = $signed(T25067) / $signed(22'h100000);
  assign T25067 = $signed(31'h21bda170) * $signed(16'h1);
  assign T25068 = T18725[1'h0:1'h0];
  assign T25069 = T18725[1'h1:1'h1];
  assign T25070 = T25091 ? T25081 : T25071;
  assign T25071 = T25080 ? twiddle4_1_333_real : twiddle4_1_332_real;
  assign twiddle4_1_332_real = T25074 + T25072;
  assign T25072 = $signed(T25073) / $signed(22'h100000);
  assign T25073 = $signed(31'h367c9a7d) * $signed(16'h0);
  assign T25074 = $signed(T25075) / $signed(22'h100000);
  assign T25075 = $signed(31'h2192e09a) * $signed(16'h1);
  assign twiddle4_1_333_real = T25078 + T25076;
  assign T25076 = $signed(T25077) / $signed(22'h100000);
  assign T25077 = $signed(31'h3696e813) * $signed(16'h0);
  assign T25078 = $signed(T25079) / $signed(22'h100000);
  assign T25079 = $signed(31'h21680b0f) * $signed(16'h1);
  assign T25080 = T18725[1'h0:1'h0];
  assign T25081 = T25090 ? twiddle4_1_335_real : twiddle4_1_334_real;
  assign twiddle4_1_334_real = T25084 + T25082;
  assign T25082 = $signed(T25083) / $signed(22'h100000);
  assign T25083 = $signed(31'h36b113fd) * $signed(16'h0);
  assign T25084 = $signed(T25085) / $signed(22'h100000);
  assign T25085 = $signed(31'h213d20e8) * $signed(16'h1);
  assign twiddle4_1_335_real = T25088 + T25086;
  assign T25086 = $signed(T25087) / $signed(22'h100000);
  assign T25087 = $signed(31'h36cb1e29) * $signed(16'h0);
  assign T25088 = $signed(T25089) / $signed(22'h100000);
  assign T25089 = $signed(31'h21122240) * $signed(16'h1);
  assign T25090 = T18725[1'h0:1'h0];
  assign T25091 = T18725[1'h1:1'h1];
  assign T25092 = T18725[2'h2:2'h2];
  assign T25093 = T18725[2'h3:2'h3];
  assign T25094 = T25207 ? T25145 : T25095;
  assign T25095 = T25144 ? T25118 : T25096;
  assign T25096 = T25117 ? T25107 : T25097;
  assign T25097 = T25106 ? twiddle4_1_337_real : twiddle4_1_336_real;
  assign twiddle4_1_336_real = T25100 + T25098;
  assign T25098 = $signed(T25099) / $signed(22'h100000);
  assign T25099 = $signed(31'h36e5068a) * $signed(16'h0);
  assign T25100 = $signed(T25101) / $signed(22'h100000);
  assign T25101 = $signed(31'h20e70f32) * $signed(16'h1);
  assign twiddle4_1_337_real = T25104 + T25102;
  assign T25102 = $signed(T25103) / $signed(22'h100000);
  assign T25103 = $signed(31'h36fecd0d) * $signed(16'h0);
  assign T25104 = $signed(T25105) / $signed(22'h100000);
  assign T25105 = $signed(31'h20bbe7d8) * $signed(16'h1);
  assign T25106 = T18725[1'h0:1'h0];
  assign T25107 = T25116 ? twiddle4_1_339_real : twiddle4_1_338_real;
  assign twiddle4_1_338_real = T25110 + T25108;
  assign T25108 = $signed(T25109) / $signed(22'h100000);
  assign T25109 = $signed(31'h371871a4) * $signed(16'h0);
  assign T25110 = $signed(T25111) / $signed(22'h100000);
  assign T25111 = $signed(31'h2090ac4d) * $signed(16'h1);
  assign twiddle4_1_339_real = T25114 + T25112;
  assign T25112 = $signed(T25113) / $signed(22'h100000);
  assign T25113 = $signed(31'h3731f43f) * $signed(16'h0);
  assign T25114 = $signed(T25115) / $signed(22'h100000);
  assign T25115 = $signed(31'h20655cab) * $signed(16'h1);
  assign T25116 = T18725[1'h0:1'h0];
  assign T25117 = T18725[1'h1:1'h1];
  assign T25118 = T25143 ? T25129 : T25119;
  assign T25119 = T25128 ? twiddle4_1_341_real : twiddle4_1_340_real;
  assign twiddle4_1_340_real = T25122 + T25120;
  assign T25120 = $signed(T25121) / $signed(22'h100000);
  assign T25121 = $signed(31'h374b54ce) * $signed(16'h0);
  assign T25122 = $signed(T25123) / $signed(22'h100000);
  assign T25123 = $signed(31'h2039f90e) * $signed(16'h1);
  assign twiddle4_1_341_real = T25126 + T25124;
  assign T25124 = $signed(T25125) / $signed(22'h100000);
  assign T25125 = $signed(31'h37649341) * $signed(16'h0);
  assign T25126 = $signed(T25127) / $signed(22'h100000);
  assign T25127 = $signed(31'h200e8190) * $signed(16'h1);
  assign T25128 = T18725[1'h0:1'h0];
  assign T25129 = T25142 ? twiddle4_1_343_real : twiddle4_1_342_real;
  assign twiddle4_1_342_real = T25132 + T25130;
  assign T25130 = $signed(T25131) / $signed(22'h100000);
  assign T25131 = $signed(31'h377daf89) * $signed(16'h0);
  assign T25132 = {T25135, T25133};
  assign T25133 = $signed(T25134) / $signed(22'h100000);
  assign T25134 = $signed(30'h1fe2f64b) * $signed(16'h1);
  assign T25135 = T25133[6'h2d:6'h2d];
  assign twiddle4_1_343_real = T25138 + T25136;
  assign T25136 = $signed(T25137) / $signed(22'h100000);
  assign T25137 = $signed(31'h3796a996) * $signed(16'h0);
  assign T25138 = {T25141, T25139};
  assign T25139 = $signed(T25140) / $signed(22'h100000);
  assign T25140 = $signed(30'h1fb7575c) * $signed(16'h1);
  assign T25141 = T25139[6'h2d:6'h2d];
  assign T25142 = T18725[1'h0:1'h0];
  assign T25143 = T18725[1'h1:1'h1];
  assign T25144 = T18725[2'h2:2'h2];
  assign T25145 = T25206 ? T25176 : T25146;
  assign T25146 = T25175 ? T25161 : T25147;
  assign T25147 = T25160 ? twiddle4_1_345_real : twiddle4_1_344_real;
  assign twiddle4_1_344_real = T25150 + T25148;
  assign T25148 = $signed(T25149) / $signed(22'h100000);
  assign T25149 = $signed(31'h37af8158) * $signed(16'h0);
  assign T25150 = {T25153, T25151};
  assign T25151 = $signed(T25152) / $signed(22'h100000);
  assign T25152 = $signed(30'h1f8ba4db) * $signed(16'h1);
  assign T25153 = T25151[6'h2d:6'h2d];
  assign twiddle4_1_345_real = T25156 + T25154;
  assign T25154 = $signed(T25155) / $signed(22'h100000);
  assign T25155 = $signed(31'h37c836c2) * $signed(16'h0);
  assign T25156 = {T25159, T25157};
  assign T25157 = $signed(T25158) / $signed(22'h100000);
  assign T25158 = $signed(30'h1f5fdee6) * $signed(16'h1);
  assign T25159 = T25157[6'h2d:6'h2d];
  assign T25160 = T18725[1'h0:1'h0];
  assign T25161 = T25174 ? twiddle4_1_347_real : twiddle4_1_346_real;
  assign twiddle4_1_346_real = T25164 + T25162;
  assign T25162 = $signed(T25163) / $signed(22'h100000);
  assign T25163 = $signed(31'h37e0c9c2) * $signed(16'h0);
  assign T25164 = {T25167, T25165};
  assign T25165 = $signed(T25166) / $signed(22'h100000);
  assign T25166 = $signed(30'h1f340596) * $signed(16'h1);
  assign T25167 = T25165[6'h2d:6'h2d];
  assign twiddle4_1_347_real = T25170 + T25168;
  assign T25168 = $signed(T25169) / $signed(22'h100000);
  assign T25169 = $signed(31'h37f93a4b) * $signed(16'h0);
  assign T25170 = {T25173, T25171};
  assign T25171 = $signed(T25172) / $signed(22'h100000);
  assign T25172 = $signed(30'h1f081906) * $signed(16'h1);
  assign T25173 = T25171[6'h2d:6'h2d];
  assign T25174 = T18725[1'h0:1'h0];
  assign T25175 = T18725[1'h1:1'h1];
  assign T25176 = T25205 ? T25191 : T25177;
  assign T25177 = T25190 ? twiddle4_1_349_real : twiddle4_1_348_real;
  assign twiddle4_1_348_real = T25180 + T25178;
  assign T25178 = $signed(T25179) / $signed(22'h100000);
  assign T25179 = $signed(31'h3811884c) * $signed(16'h0);
  assign T25180 = {T25183, T25181};
  assign T25181 = $signed(T25182) / $signed(22'h100000);
  assign T25182 = $signed(30'h1edc1952) * $signed(16'h1);
  assign T25183 = T25181[6'h2d:6'h2d];
  assign twiddle4_1_349_real = T25186 + T25184;
  assign T25184 = $signed(T25185) / $signed(22'h100000);
  assign T25185 = $signed(31'h3829b3b8) * $signed(16'h0);
  assign T25186 = {T25189, T25187};
  assign T25187 = $signed(T25188) / $signed(22'h100000);
  assign T25188 = $signed(30'h1eb00695) * $signed(16'h1);
  assign T25189 = T25187[6'h2d:6'h2d];
  assign T25190 = T18725[1'h0:1'h0];
  assign T25191 = T25204 ? twiddle4_1_351_real : twiddle4_1_350_real;
  assign twiddle4_1_350_real = T25194 + T25192;
  assign T25192 = $signed(T25193) / $signed(22'h100000);
  assign T25193 = $signed(31'h3841bc7f) * $signed(16'h0);
  assign T25194 = {T25197, T25195};
  assign T25195 = $signed(T25196) / $signed(22'h100000);
  assign T25196 = $signed(30'h1e83e0ea) * $signed(16'h1);
  assign T25197 = T25195[6'h2d:6'h2d];
  assign twiddle4_1_351_real = T25200 + T25198;
  assign T25198 = $signed(T25199) / $signed(22'h100000);
  assign T25199 = $signed(31'h3859a292) * $signed(16'h0);
  assign T25200 = {T25203, T25201};
  assign T25201 = $signed(T25202) / $signed(22'h100000);
  assign T25202 = $signed(30'h1e57a86d) * $signed(16'h1);
  assign T25203 = T25201[6'h2d:6'h2d];
  assign T25204 = T18725[1'h0:1'h0];
  assign T25205 = T18725[1'h1:1'h1];
  assign T25206 = T18725[2'h2:2'h2];
  assign T25207 = T18725[2'h3:2'h3];
  assign T25208 = T18725[3'h4:3'h4];
  assign T25209 = T25462 ? T25336 : T25210;
  assign T25210 = T25335 ? T25273 : T25211;
  assign T25211 = T25272 ? T25242 : T25212;
  assign T25212 = T25241 ? T25227 : T25213;
  assign T25213 = T25226 ? twiddle4_1_353_real : twiddle4_1_352_real;
  assign twiddle4_1_352_real = T25216 + T25214;
  assign T25214 = $signed(T25215) / $signed(22'h100000);
  assign T25215 = $signed(31'h387165e3) * $signed(16'h0);
  assign T25216 = {T25219, T25217};
  assign T25217 = $signed(T25218) / $signed(22'h100000);
  assign T25218 = $signed(30'h1e2b5d38) * $signed(16'h1);
  assign T25219 = T25217[6'h2d:6'h2d];
  assign twiddle4_1_353_real = T25222 + T25220;
  assign T25220 = $signed(T25221) / $signed(22'h100000);
  assign T25221 = $signed(31'h38890662) * $signed(16'h0);
  assign T25222 = {T25225, T25223};
  assign T25223 = $signed(T25224) / $signed(22'h100000);
  assign T25224 = $signed(30'h1dfeff66) * $signed(16'h1);
  assign T25225 = T25223[6'h2d:6'h2d];
  assign T25226 = T18725[1'h0:1'h0];
  assign T25227 = T25240 ? twiddle4_1_355_real : twiddle4_1_354_real;
  assign twiddle4_1_354_real = T25230 + T25228;
  assign T25228 = $signed(T25229) / $signed(22'h100000);
  assign T25229 = $signed(31'h38a08402) * $signed(16'h0);
  assign T25230 = {T25233, T25231};
  assign T25231 = $signed(T25232) / $signed(22'h100000);
  assign T25232 = $signed(30'h1dd28f14) * $signed(16'h1);
  assign T25233 = T25231[6'h2d:6'h2d];
  assign twiddle4_1_355_real = T25236 + T25234;
  assign T25234 = $signed(T25235) / $signed(22'h100000);
  assign T25235 = $signed(31'h38b7deb3) * $signed(16'h0);
  assign T25236 = {T25239, T25237};
  assign T25237 = $signed(T25238) / $signed(22'h100000);
  assign T25238 = $signed(30'h1da60c5c) * $signed(16'h1);
  assign T25239 = T25237[6'h2d:6'h2d];
  assign T25240 = T18725[1'h0:1'h0];
  assign T25241 = T18725[1'h1:1'h1];
  assign T25242 = T25271 ? T25257 : T25243;
  assign T25243 = T25256 ? twiddle4_1_357_real : twiddle4_1_356_real;
  assign twiddle4_1_356_real = T25246 + T25244;
  assign T25244 = $signed(T25245) / $signed(22'h100000);
  assign T25245 = $signed(31'h38cf1669) * $signed(16'h0);
  assign T25246 = {T25249, T25247};
  assign T25247 = $signed(T25248) / $signed(22'h100000);
  assign T25248 = $signed(30'h1d79775b) * $signed(16'h1);
  assign T25249 = T25247[6'h2d:6'h2d];
  assign twiddle4_1_357_real = T25252 + T25250;
  assign T25250 = $signed(T25251) / $signed(22'h100000);
  assign T25251 = $signed(31'h38e62b13) * $signed(16'h0);
  assign T25252 = {T25255, T25253};
  assign T25253 = $signed(T25254) / $signed(22'h100000);
  assign T25254 = $signed(30'h1d4cd02b) * $signed(16'h1);
  assign T25255 = T25253[6'h2d:6'h2d];
  assign T25256 = T18725[1'h0:1'h0];
  assign T25257 = T25270 ? twiddle4_1_359_real : twiddle4_1_358_real;
  assign twiddle4_1_358_real = T25260 + T25258;
  assign T25258 = $signed(T25259) / $signed(22'h100000);
  assign T25259 = $signed(31'h38fd1ca4) * $signed(16'h0);
  assign T25260 = {T25263, T25261};
  assign T25261 = $signed(T25262) / $signed(22'h100000);
  assign T25262 = $signed(30'h1d2016e8) * $signed(16'h1);
  assign T25263 = T25261[6'h2d:6'h2d];
  assign twiddle4_1_359_real = T25266 + T25264;
  assign T25264 = $signed(T25265) / $signed(22'h100000);
  assign T25265 = $signed(31'h3913eb0e) * $signed(16'h0);
  assign T25266 = {T25269, T25267};
  assign T25267 = $signed(T25268) / $signed(22'h100000);
  assign T25268 = $signed(30'h1cf34bae) * $signed(16'h1);
  assign T25269 = T25267[6'h2d:6'h2d];
  assign T25270 = T18725[1'h0:1'h0];
  assign T25271 = T18725[1'h1:1'h1];
  assign T25272 = T18725[2'h2:2'h2];
  assign T25273 = T25334 ? T25304 : T25274;
  assign T25274 = T25303 ? T25289 : T25275;
  assign T25275 = T25288 ? twiddle4_1_361_real : twiddle4_1_360_real;
  assign twiddle4_1_360_real = T25278 + T25276;
  assign T25276 = $signed(T25277) / $signed(22'h100000);
  assign T25277 = $signed(31'h392a9642) * $signed(16'h0);
  assign T25278 = {T25281, T25279};
  assign T25279 = $signed(T25280) / $signed(22'h100000);
  assign T25280 = $signed(30'h1cc66e99) * $signed(16'h1);
  assign T25281 = T25279[6'h2d:6'h2d];
  assign twiddle4_1_361_real = T25284 + T25282;
  assign T25282 = $signed(T25283) / $signed(22'h100000);
  assign T25283 = $signed(31'h39411e33) * $signed(16'h0);
  assign T25284 = {T25287, T25285};
  assign T25285 = $signed(T25286) / $signed(22'h100000);
  assign T25286 = $signed(30'h1c997fc3) * $signed(16'h1);
  assign T25287 = T25285[6'h2d:6'h2d];
  assign T25288 = T18725[1'h0:1'h0];
  assign T25289 = T25302 ? twiddle4_1_363_real : twiddle4_1_362_real;
  assign twiddle4_1_362_real = T25292 + T25290;
  assign T25290 = $signed(T25291) / $signed(22'h100000);
  assign T25291 = $signed(31'h395782d3) * $signed(16'h0);
  assign T25292 = {T25295, T25293};
  assign T25293 = $signed(T25294) / $signed(22'h100000);
  assign T25294 = $signed(30'h1c6c7f49) * $signed(16'h1);
  assign T25295 = T25293[6'h2d:6'h2d];
  assign twiddle4_1_363_real = T25298 + T25296;
  assign T25296 = $signed(T25297) / $signed(22'h100000);
  assign T25297 = $signed(31'h396dc414) * $signed(16'h0);
  assign T25298 = {T25301, T25299};
  assign T25299 = $signed(T25300) / $signed(22'h100000);
  assign T25300 = $signed(30'h1c3f6d47) * $signed(16'h1);
  assign T25301 = T25299[6'h2d:6'h2d];
  assign T25302 = T18725[1'h0:1'h0];
  assign T25303 = T18725[1'h1:1'h1];
  assign T25304 = T25333 ? T25319 : T25305;
  assign T25305 = T25318 ? twiddle4_1_365_real : twiddle4_1_364_real;
  assign twiddle4_1_364_real = T25308 + T25306;
  assign T25306 = $signed(T25307) / $signed(22'h100000);
  assign T25307 = $signed(31'h3983e1e7) * $signed(16'h0);
  assign T25308 = {T25311, T25309};
  assign T25309 = $signed(T25310) / $signed(22'h100000);
  assign T25310 = $signed(30'h1c1249d8) * $signed(16'h1);
  assign T25311 = T25309[6'h2d:6'h2d];
  assign twiddle4_1_365_real = T25314 + T25312;
  assign T25312 = $signed(T25313) / $signed(22'h100000);
  assign T25313 = $signed(31'h3999dc41) * $signed(16'h0);
  assign T25314 = {T25317, T25315};
  assign T25315 = $signed(T25316) / $signed(22'h100000);
  assign T25316 = $signed(30'h1be51517) * $signed(16'h1);
  assign T25317 = T25315[6'h2d:6'h2d];
  assign T25318 = T18725[1'h0:1'h0];
  assign T25319 = T25332 ? twiddle4_1_367_real : twiddle4_1_366_real;
  assign twiddle4_1_366_real = T25322 + T25320;
  assign T25320 = $signed(T25321) / $signed(22'h100000);
  assign T25321 = $signed(31'h39afb313) * $signed(16'h0);
  assign T25322 = {T25325, T25323};
  assign T25323 = $signed(T25324) / $signed(22'h100000);
  assign T25324 = $signed(30'h1bb7cf23) * $signed(16'h1);
  assign T25325 = T25323[6'h2d:6'h2d];
  assign twiddle4_1_367_real = T25328 + T25326;
  assign T25326 = $signed(T25327) / $signed(22'h100000);
  assign T25327 = $signed(31'h39c5664f) * $signed(16'h0);
  assign T25328 = {T25331, T25329};
  assign T25329 = $signed(T25330) / $signed(22'h100000);
  assign T25330 = $signed(30'h1b8a7814) * $signed(16'h1);
  assign T25331 = T25329[6'h2d:6'h2d];
  assign T25332 = T18725[1'h0:1'h0];
  assign T25333 = T18725[1'h1:1'h1];
  assign T25334 = T18725[2'h2:2'h2];
  assign T25335 = T18725[2'h3:2'h3];
  assign T25336 = T25461 ? T25399 : T25337;
  assign T25337 = T25398 ? T25368 : T25338;
  assign T25338 = T25367 ? T25353 : T25339;
  assign T25339 = T25352 ? twiddle4_1_369_real : twiddle4_1_368_real;
  assign twiddle4_1_368_real = T25342 + T25340;
  assign T25340 = $signed(T25341) / $signed(22'h100000);
  assign T25341 = $signed(31'h39daf5e8) * $signed(16'h0);
  assign T25342 = {T25345, T25343};
  assign T25343 = $signed(T25344) / $signed(22'h100000);
  assign T25344 = $signed(30'h1b5d1009) * $signed(16'h1);
  assign T25345 = T25343[6'h2d:6'h2d];
  assign twiddle4_1_369_real = T25348 + T25346;
  assign T25346 = $signed(T25347) / $signed(22'h100000);
  assign T25347 = $signed(31'h39f061d1) * $signed(16'h0);
  assign T25348 = {T25351, T25349};
  assign T25349 = $signed(T25350) / $signed(22'h100000);
  assign T25350 = $signed(30'h1b2f971d) * $signed(16'h1);
  assign T25351 = T25349[6'h2d:6'h2d];
  assign T25352 = T18725[1'h0:1'h0];
  assign T25353 = T25366 ? twiddle4_1_371_real : twiddle4_1_370_real;
  assign twiddle4_1_370_real = T25356 + T25354;
  assign T25354 = $signed(T25355) / $signed(22'h100000);
  assign T25355 = $signed(31'h3a05a9fd) * $signed(16'h0);
  assign T25356 = {T25359, T25357};
  assign T25357 = $signed(T25358) / $signed(22'h100000);
  assign T25358 = $signed(30'h1b020d6c) * $signed(16'h1);
  assign T25359 = T25357[6'h2d:6'h2d];
  assign twiddle4_1_371_real = T25362 + T25360;
  assign T25360 = $signed(T25361) / $signed(22'h100000);
  assign T25361 = $signed(31'h3a1ace5e) * $signed(16'h0);
  assign T25362 = {T25365, T25363};
  assign T25363 = $signed(T25364) / $signed(22'h100000);
  assign T25364 = $signed(30'h1ad47312) * $signed(16'h1);
  assign T25365 = T25363[6'h2d:6'h2d];
  assign T25366 = T18725[1'h0:1'h0];
  assign T25367 = T18725[1'h1:1'h1];
  assign T25368 = T25397 ? T25383 : T25369;
  assign T25369 = T25382 ? twiddle4_1_373_real : twiddle4_1_372_real;
  assign twiddle4_1_372_real = T25372 + T25370;
  assign T25370 = $signed(T25371) / $signed(22'h100000);
  assign T25371 = $signed(31'h3a2fcee8) * $signed(16'h0);
  assign T25372 = {T25375, T25373};
  assign T25373 = $signed(T25374) / $signed(22'h100000);
  assign T25374 = $signed(30'h1aa6c82b) * $signed(16'h1);
  assign T25375 = T25373[6'h2d:6'h2d];
  assign twiddle4_1_373_real = T25378 + T25376;
  assign T25376 = $signed(T25377) / $signed(22'h100000);
  assign T25377 = $signed(31'h3a44ab8d) * $signed(16'h0);
  assign T25378 = {T25381, T25379};
  assign T25379 = $signed(T25380) / $signed(22'h100000);
  assign T25380 = $signed(30'h1a790cd3) * $signed(16'h1);
  assign T25381 = T25379[6'h2d:6'h2d];
  assign T25382 = T18725[1'h0:1'h0];
  assign T25383 = T25396 ? twiddle4_1_375_real : twiddle4_1_374_real;
  assign twiddle4_1_374_real = T25386 + T25384;
  assign T25384 = $signed(T25385) / $signed(22'h100000);
  assign T25385 = $signed(31'h3a596441) * $signed(16'h0);
  assign T25386 = {T25389, T25387};
  assign T25387 = $signed(T25388) / $signed(22'h100000);
  assign T25388 = $signed(30'h1a4b4127) * $signed(16'h1);
  assign T25389 = T25387[6'h2d:6'h2d];
  assign twiddle4_1_375_real = T25392 + T25390;
  assign T25390 = $signed(T25391) / $signed(22'h100000);
  assign T25391 = $signed(31'h3a6df8f7) * $signed(16'h0);
  assign T25392 = {T25395, T25393};
  assign T25393 = $signed(T25394) / $signed(22'h100000);
  assign T25394 = $signed(30'h1a1d6543) * $signed(16'h1);
  assign T25395 = T25393[6'h2d:6'h2d];
  assign T25396 = T18725[1'h0:1'h0];
  assign T25397 = T18725[1'h1:1'h1];
  assign T25398 = T18725[2'h2:2'h2];
  assign T25399 = T25460 ? T25430 : T25400;
  assign T25400 = T25429 ? T25415 : T25401;
  assign T25401 = T25414 ? twiddle4_1_377_real : twiddle4_1_376_real;
  assign twiddle4_1_376_real = T25404 + T25402;
  assign T25402 = $signed(T25403) / $signed(22'h100000);
  assign T25403 = $signed(31'h3a8269a2) * $signed(16'h0);
  assign T25404 = {T25407, T25405};
  assign T25405 = $signed(T25406) / $signed(22'h100000);
  assign T25406 = $signed(30'h19ef7943) * $signed(16'h1);
  assign T25407 = T25405[6'h2d:6'h2d];
  assign twiddle4_1_377_real = T25410 + T25408;
  assign T25408 = $signed(T25409) / $signed(22'h100000);
  assign T25409 = $signed(31'h3a96b636) * $signed(16'h0);
  assign T25410 = {T25413, T25411};
  assign T25411 = $signed(T25412) / $signed(22'h100000);
  assign T25412 = $signed(30'h19c17d44) * $signed(16'h1);
  assign T25413 = T25411[6'h2d:6'h2d];
  assign T25414 = T18725[1'h0:1'h0];
  assign T25415 = T25428 ? twiddle4_1_379_real : twiddle4_1_378_real;
  assign twiddle4_1_378_real = T25418 + T25416;
  assign T25416 = $signed(T25417) / $signed(22'h100000);
  assign T25417 = $signed(31'h3aaadea5) * $signed(16'h0);
  assign T25418 = {T25421, T25419};
  assign T25419 = $signed(T25420) / $signed(22'h100000);
  assign T25420 = $signed(30'h19937161) * $signed(16'h1);
  assign T25421 = T25419[6'h2d:6'h2d];
  assign twiddle4_1_379_real = T25424 + T25422;
  assign T25422 = $signed(T25423) / $signed(22'h100000);
  assign T25423 = $signed(31'h3abee2e5) * $signed(16'h0);
  assign T25424 = {T25427, T25425};
  assign T25425 = $signed(T25426) / $signed(22'h100000);
  assign T25426 = $signed(30'h196555b7) * $signed(16'h1);
  assign T25427 = T25425[6'h2d:6'h2d];
  assign T25428 = T18725[1'h0:1'h0];
  assign T25429 = T18725[1'h1:1'h1];
  assign T25430 = T25459 ? T25445 : T25431;
  assign T25431 = T25444 ? twiddle4_1_381_real : twiddle4_1_380_real;
  assign twiddle4_1_380_real = T25434 + T25432;
  assign T25432 = $signed(T25433) / $signed(22'h100000);
  assign T25433 = $signed(31'h3ad2c2e7) * $signed(16'h0);
  assign T25434 = {T25437, T25435};
  assign T25435 = $signed(T25436) / $signed(22'h100000);
  assign T25436 = $signed(30'h19372a63) * $signed(16'h1);
  assign T25437 = T25435[6'h2d:6'h2d];
  assign twiddle4_1_381_real = T25440 + T25438;
  assign T25438 = $signed(T25439) / $signed(22'h100000);
  assign T25439 = $signed(31'h3ae67ea1) * $signed(16'h0);
  assign T25440 = {T25443, T25441};
  assign T25441 = $signed(T25442) / $signed(22'h100000);
  assign T25442 = $signed(30'h1908ef81) * $signed(16'h1);
  assign T25443 = T25441[6'h2d:6'h2d];
  assign T25444 = T18725[1'h0:1'h0];
  assign T25445 = T25458 ? twiddle4_1_383_real : twiddle4_1_382_real;
  assign twiddle4_1_382_real = T25448 + T25446;
  assign T25446 = $signed(T25447) / $signed(22'h100000);
  assign T25447 = $signed(31'h3afa1605) * $signed(16'h0);
  assign T25448 = {T25451, T25449};
  assign T25449 = $signed(T25450) / $signed(22'h100000);
  assign T25450 = $signed(30'h18daa52e) * $signed(16'h1);
  assign T25451 = T25449[6'h2d:6'h2d];
  assign twiddle4_1_383_real = T25454 + T25452;
  assign T25452 = $signed(T25453) / $signed(22'h100000);
  assign T25453 = $signed(31'h3b0d8908) * $signed(16'h0);
  assign T25454 = {T25457, T25455};
  assign T25455 = $signed(T25456) / $signed(22'h100000);
  assign T25456 = $signed(30'h18ac4b86) * $signed(16'h1);
  assign T25457 = T25455[6'h2d:6'h2d];
  assign T25458 = T18725[1'h0:1'h0];
  assign T25459 = T18725[1'h1:1'h1];
  assign T25460 = T18725[2'h2:2'h2];
  assign T25461 = T18725[2'h3:2'h3];
  assign T25462 = T18725[3'h4:3'h4];
  assign T25463 = T18725[3'h5:3'h5];
  assign T25464 = T18725[3'h6:3'h6];
  assign T25465 = T26568 ? T25994 : T25466;
  assign T25466 = T25993 ? T25721 : T25467;
  assign T25467 = T25720 ? T25594 : T25468;
  assign T25468 = T25593 ? T25531 : T25469;
  assign T25469 = T25530 ? T25500 : T25470;
  assign T25470 = T25499 ? T25485 : T25471;
  assign T25471 = T25484 ? twiddle4_1_385_real : twiddle4_1_384_real;
  assign twiddle4_1_384_real = T25474 + T25472;
  assign T25472 = $signed(T25473) / $signed(22'h100000);
  assign T25473 = $signed(31'h3b20d79e) * $signed(16'h0);
  assign T25474 = {T25477, T25475};
  assign T25475 = $signed(T25476) / $signed(22'h100000);
  assign T25476 = $signed(30'h187de2a6) * $signed(16'h1);
  assign T25477 = T25475[6'h2d:6'h2d];
  assign twiddle4_1_385_real = T25480 + T25478;
  assign T25478 = $signed(T25479) / $signed(22'h100000);
  assign T25479 = $signed(31'h3b3401bb) * $signed(16'h0);
  assign T25480 = {T25483, T25481};
  assign T25481 = $signed(T25482) / $signed(22'h100000);
  assign T25482 = $signed(30'h184f6aaa) * $signed(16'h1);
  assign T25483 = T25481[6'h2d:6'h2d];
  assign T25484 = T18725[1'h0:1'h0];
  assign T25485 = T25498 ? twiddle4_1_387_real : twiddle4_1_386_real;
  assign twiddle4_1_386_real = T25488 + T25486;
  assign T25486 = $signed(T25487) / $signed(22'h100000);
  assign T25487 = $signed(31'h3b470752) * $signed(16'h0);
  assign T25488 = {T25491, T25489};
  assign T25489 = $signed(T25490) / $signed(22'h100000);
  assign T25490 = $signed(30'h1820e3b0) * $signed(16'h1);
  assign T25491 = T25489[6'h2d:6'h2d];
  assign twiddle4_1_387_real = T25494 + T25492;
  assign T25492 = $signed(T25493) / $signed(22'h100000);
  assign T25493 = $signed(31'h3b59e859) * $signed(16'h0);
  assign T25494 = {T25497, T25495};
  assign T25495 = $signed(T25496) / $signed(22'h100000);
  assign T25496 = $signed(30'h17f24dd3) * $signed(16'h1);
  assign T25497 = T25495[6'h2d:6'h2d];
  assign T25498 = T18725[1'h0:1'h0];
  assign T25499 = T18725[1'h1:1'h1];
  assign T25500 = T25529 ? T25515 : T25501;
  assign T25501 = T25514 ? twiddle4_1_389_real : twiddle4_1_388_real;
  assign twiddle4_1_388_real = T25504 + T25502;
  assign T25502 = $signed(T25503) / $signed(22'h100000);
  assign T25503 = $signed(31'h3b6ca4c4) * $signed(16'h0);
  assign T25504 = {T25507, T25505};
  assign T25505 = $signed(T25506) / $signed(22'h100000);
  assign T25506 = $signed(30'h17c3a931) * $signed(16'h1);
  assign T25507 = T25505[6'h2d:6'h2d];
  assign twiddle4_1_389_real = T25510 + T25508;
  assign T25508 = $signed(T25509) / $signed(22'h100000);
  assign T25509 = $signed(31'h3b7f3c87) * $signed(16'h0);
  assign T25510 = {T25513, T25511};
  assign T25511 = $signed(T25512) / $signed(22'h100000);
  assign T25512 = $signed(30'h1794f5e6) * $signed(16'h1);
  assign T25513 = T25511[6'h2d:6'h2d];
  assign T25514 = T18725[1'h0:1'h0];
  assign T25515 = T25528 ? twiddle4_1_391_real : twiddle4_1_390_real;
  assign twiddle4_1_390_real = T25518 + T25516;
  assign T25516 = $signed(T25517) / $signed(22'h100000);
  assign T25517 = $signed(31'h3b91af96) * $signed(16'h0);
  assign T25518 = {T25521, T25519};
  assign T25519 = $signed(T25520) / $signed(22'h100000);
  assign T25520 = $signed(30'h1766340f) * $signed(16'h1);
  assign T25521 = T25519[6'h2d:6'h2d];
  assign twiddle4_1_391_real = T25524 + T25522;
  assign T25522 = $signed(T25523) / $signed(22'h100000);
  assign T25523 = $signed(31'h3ba3fde7) * $signed(16'h0);
  assign T25524 = {T25527, T25525};
  assign T25525 = $signed(T25526) / $signed(22'h100000);
  assign T25526 = $signed(30'h173763c9) * $signed(16'h1);
  assign T25527 = T25525[6'h2d:6'h2d];
  assign T25528 = T18725[1'h0:1'h0];
  assign T25529 = T18725[1'h1:1'h1];
  assign T25530 = T18725[2'h2:2'h2];
  assign T25531 = T25592 ? T25562 : T25532;
  assign T25532 = T25561 ? T25547 : T25533;
  assign T25533 = T25546 ? twiddle4_1_393_real : twiddle4_1_392_real;
  assign twiddle4_1_392_real = T25536 + T25534;
  assign T25534 = $signed(T25535) / $signed(22'h100000);
  assign T25535 = $signed(31'h3bb6276d) * $signed(16'h0);
  assign T25536 = {T25539, T25537};
  assign T25537 = $signed(T25538) / $signed(22'h100000);
  assign T25538 = $signed(30'h17088530) * $signed(16'h1);
  assign T25539 = T25537[6'h2d:6'h2d];
  assign twiddle4_1_393_real = T25542 + T25540;
  assign T25540 = $signed(T25541) / $signed(22'h100000);
  assign T25541 = $signed(31'h3bc82c1e) * $signed(16'h0);
  assign T25542 = {T25545, T25543};
  assign T25543 = $signed(T25544) / $signed(22'h100000);
  assign T25544 = $signed(30'h16d99863) * $signed(16'h1);
  assign T25545 = T25543[6'h2d:6'h2d];
  assign T25546 = T18725[1'h0:1'h0];
  assign T25547 = T25560 ? twiddle4_1_395_real : twiddle4_1_394_real;
  assign twiddle4_1_394_real = T25550 + T25548;
  assign T25548 = $signed(T25549) / $signed(22'h100000);
  assign T25549 = $signed(31'h3bda0bef) * $signed(16'h0);
  assign T25550 = {T25553, T25551};
  assign T25551 = $signed(T25552) / $signed(22'h100000);
  assign T25552 = $signed(30'h16aa9d7d) * $signed(16'h1);
  assign T25553 = T25551[6'h2d:6'h2d];
  assign twiddle4_1_395_real = T25556 + T25554;
  assign T25554 = $signed(T25555) / $signed(22'h100000);
  assign T25555 = $signed(31'h3bebc6d5) * $signed(16'h0);
  assign T25556 = {T25559, T25557};
  assign T25557 = $signed(T25558) / $signed(22'h100000);
  assign T25558 = $signed(30'h167b949c) * $signed(16'h1);
  assign T25559 = T25557[6'h2d:6'h2d];
  assign T25560 = T18725[1'h0:1'h0];
  assign T25561 = T18725[1'h1:1'h1];
  assign T25562 = T25591 ? T25577 : T25563;
  assign T25563 = T25576 ? twiddle4_1_397_real : twiddle4_1_396_real;
  assign twiddle4_1_396_real = T25566 + T25564;
  assign T25564 = $signed(T25565) / $signed(22'h100000);
  assign T25565 = $signed(31'h3bfd5cc4) * $signed(16'h0);
  assign T25566 = {T25569, T25567};
  assign T25567 = $signed(T25568) / $signed(22'h100000);
  assign T25568 = $signed(30'h164c7ddd) * $signed(16'h1);
  assign T25569 = T25567[6'h2d:6'h2d];
  assign twiddle4_1_397_real = T25572 + T25570;
  assign T25570 = $signed(T25571) / $signed(22'h100000);
  assign T25571 = $signed(31'h3c0ecdb2) * $signed(16'h0);
  assign T25572 = {T25575, T25573};
  assign T25573 = $signed(T25574) / $signed(22'h100000);
  assign T25574 = $signed(30'h161d595c) * $signed(16'h1);
  assign T25575 = T25573[6'h2d:6'h2d];
  assign T25576 = T18725[1'h0:1'h0];
  assign T25577 = T25590 ? twiddle4_1_399_real : twiddle4_1_398_real;
  assign twiddle4_1_398_real = T25580 + T25578;
  assign T25578 = $signed(T25579) / $signed(22'h100000);
  assign T25579 = $signed(31'h3c201994) * $signed(16'h0);
  assign T25580 = {T25583, T25581};
  assign T25581 = $signed(T25582) / $signed(22'h100000);
  assign T25582 = $signed(30'h15ee2737) * $signed(16'h1);
  assign T25583 = T25581[6'h2d:6'h2d];
  assign twiddle4_1_399_real = T25586 + T25584;
  assign T25584 = $signed(T25585) / $signed(22'h100000);
  assign T25585 = $signed(31'h3c31405f) * $signed(16'h0);
  assign T25586 = {T25589, T25587};
  assign T25587 = $signed(T25588) / $signed(22'h100000);
  assign T25588 = $signed(30'h15bee78b) * $signed(16'h1);
  assign T25589 = T25587[6'h2d:6'h2d];
  assign T25590 = T18725[1'h0:1'h0];
  assign T25591 = T18725[1'h1:1'h1];
  assign T25592 = T18725[2'h2:2'h2];
  assign T25593 = T18725[2'h3:2'h3];
  assign T25594 = T25719 ? T25657 : T25595;
  assign T25595 = T25656 ? T25626 : T25596;
  assign T25596 = T25625 ? T25611 : T25597;
  assign T25597 = T25610 ? twiddle4_1_401_real : twiddle4_1_400_real;
  assign twiddle4_1_400_real = T25600 + T25598;
  assign T25598 = $signed(T25599) / $signed(22'h100000);
  assign T25599 = $signed(31'h3c424209) * $signed(16'h0);
  assign T25600 = {T25603, T25601};
  assign T25601 = $signed(T25602) / $signed(22'h100000);
  assign T25602 = $signed(30'h158f9a75) * $signed(16'h1);
  assign T25603 = T25601[6'h2d:6'h2d];
  assign twiddle4_1_401_real = T25606 + T25604;
  assign T25604 = $signed(T25605) / $signed(22'h100000);
  assign T25605 = $signed(31'h3c531e88) * $signed(16'h0);
  assign T25606 = {T25609, T25607};
  assign T25607 = $signed(T25608) / $signed(22'h100000);
  assign T25608 = $signed(30'h15604012) * $signed(16'h1);
  assign T25609 = T25607[6'h2d:6'h2d];
  assign T25610 = T18725[1'h0:1'h0];
  assign T25611 = T25624 ? twiddle4_1_403_real : twiddle4_1_402_real;
  assign twiddle4_1_402_real = T25614 + T25612;
  assign T25612 = $signed(T25613) / $signed(22'h100000);
  assign T25613 = $signed(31'h3c63d5d0) * $signed(16'h0);
  assign T25614 = {T25617, T25615};
  assign T25615 = $signed(T25616) / $signed(22'h100000);
  assign T25616 = $signed(30'h1530d880) * $signed(16'h1);
  assign T25617 = T25615[6'h2d:6'h2d];
  assign twiddle4_1_403_real = T25620 + T25618;
  assign T25618 = $signed(T25619) / $signed(22'h100000);
  assign T25619 = $signed(31'h3c7467d8) * $signed(16'h0);
  assign T25620 = {T25623, T25621};
  assign T25621 = $signed(T25622) / $signed(22'h100000);
  assign T25622 = $signed(30'h150163dc) * $signed(16'h1);
  assign T25623 = T25621[6'h2d:6'h2d];
  assign T25624 = T18725[1'h0:1'h0];
  assign T25625 = T18725[1'h1:1'h1];
  assign T25626 = T25655 ? T25641 : T25627;
  assign T25627 = T25640 ? twiddle4_1_405_real : twiddle4_1_404_real;
  assign twiddle4_1_404_real = T25630 + T25628;
  assign T25628 = $signed(T25629) / $signed(22'h100000);
  assign T25629 = $signed(31'h3c84d496) * $signed(16'h0);
  assign T25630 = {T25633, T25631};
  assign T25631 = $signed(T25632) / $signed(22'h100000);
  assign T25632 = $signed(30'h14d1e242) * $signed(16'h1);
  assign T25633 = T25631[6'h2d:6'h2d];
  assign twiddle4_1_405_real = T25636 + T25634;
  assign T25634 = $signed(T25635) / $signed(22'h100000);
  assign T25635 = $signed(31'h3c951bff) * $signed(16'h0);
  assign T25636 = {T25639, T25637};
  assign T25637 = $signed(T25638) / $signed(22'h100000);
  assign T25638 = $signed(30'h14a253d1) * $signed(16'h1);
  assign T25639 = T25637[6'h2d:6'h2d];
  assign T25640 = T18725[1'h0:1'h0];
  assign T25641 = T25654 ? twiddle4_1_407_real : twiddle4_1_406_real;
  assign twiddle4_1_406_real = T25644 + T25642;
  assign T25642 = $signed(T25643) / $signed(22'h100000);
  assign T25643 = $signed(31'h3ca53e08) * $signed(16'h0);
  assign T25644 = {T25647, T25645};
  assign T25645 = $signed(T25646) / $signed(22'h100000);
  assign T25646 = $signed(30'h1472b8a5) * $signed(16'h1);
  assign T25647 = T25645[6'h2d:6'h2d];
  assign twiddle4_1_407_real = T25650 + T25648;
  assign T25648 = $signed(T25649) / $signed(22'h100000);
  assign T25649 = $signed(31'h3cb53aaa) * $signed(16'h0);
  assign T25650 = {T25653, T25651};
  assign T25651 = $signed(T25652) / $signed(22'h100000);
  assign T25652 = $signed(30'h144310dc) * $signed(16'h1);
  assign T25653 = T25651[6'h2d:6'h2d];
  assign T25654 = T18725[1'h0:1'h0];
  assign T25655 = T18725[1'h1:1'h1];
  assign T25656 = T18725[2'h2:2'h2];
  assign T25657 = T25718 ? T25688 : T25658;
  assign T25658 = T25687 ? T25673 : T25659;
  assign T25659 = T25672 ? twiddle4_1_409_real : twiddle4_1_408_real;
  assign twiddle4_1_408_real = T25662 + T25660;
  assign T25660 = $signed(T25661) / $signed(22'h100000);
  assign T25661 = $signed(31'h3cc511d8) * $signed(16'h0);
  assign T25662 = {T25665, T25663};
  assign T25663 = $signed(T25664) / $signed(22'h100000);
  assign T25664 = $signed(30'h14135c94) * $signed(16'h1);
  assign T25665 = T25663[6'h2d:6'h2d];
  assign twiddle4_1_409_real = T25668 + T25666;
  assign T25666 = $signed(T25667) / $signed(22'h100000);
  assign T25667 = $signed(31'h3cd4c38a) * $signed(16'h0);
  assign T25668 = {T25671, T25669};
  assign T25669 = $signed(T25670) / $signed(22'h100000);
  assign T25670 = $signed(30'h13e39be9) * $signed(16'h1);
  assign T25671 = T25669[6'h2d:6'h2d];
  assign T25672 = T18725[1'h0:1'h0];
  assign T25673 = T25686 ? twiddle4_1_411_real : twiddle4_1_410_real;
  assign twiddle4_1_410_real = T25676 + T25674;
  assign T25674 = $signed(T25675) / $signed(22'h100000);
  assign T25675 = $signed(31'h3ce44fb6) * $signed(16'h0);
  assign T25676 = {T25679, T25677};
  assign T25677 = $signed(T25678) / $signed(22'h100000);
  assign T25678 = $signed(30'h13b3cefa) * $signed(16'h1);
  assign T25679 = T25677[6'h2d:6'h2d];
  assign twiddle4_1_411_real = T25682 + T25680;
  assign T25680 = $signed(T25681) / $signed(22'h100000);
  assign T25681 = $signed(31'h3cf3b653) * $signed(16'h0);
  assign T25682 = {T25685, T25683};
  assign T25683 = $signed(T25684) / $signed(22'h100000);
  assign T25684 = $signed(30'h1383f5e3) * $signed(16'h1);
  assign T25685 = T25683[6'h2d:6'h2d];
  assign T25686 = T18725[1'h0:1'h0];
  assign T25687 = T18725[1'h1:1'h1];
  assign T25688 = T25717 ? T25703 : T25689;
  assign T25689 = T25702 ? twiddle4_1_413_real : twiddle4_1_412_real;
  assign twiddle4_1_412_real = T25692 + T25690;
  assign T25690 = $signed(T25691) / $signed(22'h100000);
  assign T25691 = $signed(31'h3d02f756) * $signed(16'h0);
  assign T25692 = {T25695, T25693};
  assign T25693 = $signed(T25694) / $signed(22'h100000);
  assign T25694 = $signed(30'h135410c2) * $signed(16'h1);
  assign T25695 = T25693[6'h2d:6'h2d];
  assign twiddle4_1_413_real = T25698 + T25696;
  assign T25696 = $signed(T25697) / $signed(22'h100000);
  assign T25697 = $signed(31'h3d1212b7) * $signed(16'h0);
  assign T25698 = {T25701, T25699};
  assign T25699 = $signed(T25700) / $signed(22'h100000);
  assign T25700 = $signed(30'h13241fb6) * $signed(16'h1);
  assign T25701 = T25699[6'h2d:6'h2d];
  assign T25702 = T18725[1'h0:1'h0];
  assign T25703 = T25716 ? twiddle4_1_415_real : twiddle4_1_414_real;
  assign twiddle4_1_414_real = T25706 + T25704;
  assign T25704 = $signed(T25705) / $signed(22'h100000);
  assign T25705 = $signed(31'h3d21086c) * $signed(16'h0);
  assign T25706 = {T25709, T25707};
  assign T25707 = $signed(T25708) / $signed(22'h100000);
  assign T25708 = $signed(30'h12f422da) * $signed(16'h1);
  assign T25709 = T25707[6'h2d:6'h2d];
  assign twiddle4_1_415_real = T25712 + T25710;
  assign T25710 = $signed(T25711) / $signed(22'h100000);
  assign T25711 = $signed(31'h3d2fd86c) * $signed(16'h0);
  assign T25712 = {T25715, T25713};
  assign T25713 = $signed(T25714) / $signed(22'h100000);
  assign T25714 = $signed(30'h12c41a4e) * $signed(16'h1);
  assign T25715 = T25713[6'h2d:6'h2d];
  assign T25716 = T18725[1'h0:1'h0];
  assign T25717 = T18725[1'h1:1'h1];
  assign T25718 = T18725[2'h2:2'h2];
  assign T25719 = T18725[2'h3:2'h3];
  assign T25720 = T18725[3'h4:3'h4];
  assign T25721 = T25992 ? T25850 : T25722;
  assign T25722 = T25849 ? T25785 : T25723;
  assign T25723 = T25784 ? T25754 : T25724;
  assign T25724 = T25753 ? T25739 : T25725;
  assign T25725 = T25738 ? twiddle4_1_417_real : twiddle4_1_416_real;
  assign twiddle4_1_416_real = T25728 + T25726;
  assign T25726 = $signed(T25727) / $signed(22'h100000);
  assign T25727 = $signed(31'h3d3e82ad) * $signed(16'h0);
  assign T25728 = {T25731, T25729};
  assign T25729 = $signed(T25730) / $signed(22'h100000);
  assign T25730 = $signed(30'h1294062e) * $signed(16'h1);
  assign T25731 = T25729[6'h2d:6'h2d];
  assign twiddle4_1_417_real = T25734 + T25732;
  assign T25732 = $signed(T25733) / $signed(22'h100000);
  assign T25733 = $signed(31'h3d4d0727) * $signed(16'h0);
  assign T25734 = {T25737, T25735};
  assign T25735 = $signed(T25736) / $signed(22'h100000);
  assign T25736 = $signed(30'h1263e699) * $signed(16'h1);
  assign T25737 = T25735[6'h2d:6'h2d];
  assign T25738 = T18725[1'h0:1'h0];
  assign T25739 = T25752 ? twiddle4_1_419_real : twiddle4_1_418_real;
  assign twiddle4_1_418_real = T25742 + T25740;
  assign T25740 = $signed(T25741) / $signed(22'h100000);
  assign T25741 = $signed(31'h3d5b65d1) * $signed(16'h0);
  assign T25742 = {T25745, T25743};
  assign T25743 = $signed(T25744) / $signed(22'h100000);
  assign T25744 = $signed(30'h1233bbab) * $signed(16'h1);
  assign T25745 = T25743[6'h2d:6'h2d];
  assign twiddle4_1_419_real = T25748 + T25746;
  assign T25746 = $signed(T25747) / $signed(22'h100000);
  assign T25747 = $signed(31'h3d699ea2) * $signed(16'h0);
  assign T25748 = {T25751, T25749};
  assign T25749 = $signed(T25750) / $signed(22'h100000);
  assign T25750 = $signed(30'h12038583) * $signed(16'h1);
  assign T25751 = T25749[6'h2d:6'h2d];
  assign T25752 = T18725[1'h0:1'h0];
  assign T25753 = T18725[1'h1:1'h1];
  assign T25754 = T25783 ? T25769 : T25755;
  assign T25755 = T25768 ? twiddle4_1_421_real : twiddle4_1_420_real;
  assign twiddle4_1_420_real = T25758 + T25756;
  assign T25756 = $signed(T25757) / $signed(22'h100000);
  assign T25757 = $signed(31'h3d77b191) * $signed(16'h0);
  assign T25758 = {T25761, T25759};
  assign T25759 = $signed(T25760) / $signed(22'h100000);
  assign T25760 = $signed(30'h11d3443f) * $signed(16'h1);
  assign T25761 = T25759[6'h2d:6'h2d];
  assign twiddle4_1_421_real = T25764 + T25762;
  assign T25762 = $signed(T25763) / $signed(22'h100000);
  assign T25763 = $signed(31'h3d859e96) * $signed(16'h0);
  assign T25764 = {T25767, T25765};
  assign T25765 = $signed(T25766) / $signed(22'h100000);
  assign T25766 = $signed(30'h11a2f7fb) * $signed(16'h1);
  assign T25767 = T25765[6'h2d:6'h2d];
  assign T25768 = T18725[1'h0:1'h0];
  assign T25769 = T25782 ? twiddle4_1_423_real : twiddle4_1_422_real;
  assign twiddle4_1_422_real = T25772 + T25770;
  assign T25770 = $signed(T25771) / $signed(22'h100000);
  assign T25771 = $signed(31'h3d9365a7) * $signed(16'h0);
  assign T25772 = {T25775, T25773};
  assign T25773 = $signed(T25774) / $signed(22'h100000);
  assign T25774 = $signed(30'h1172a0d7) * $signed(16'h1);
  assign T25775 = T25773[6'h2d:6'h2d];
  assign twiddle4_1_423_real = T25778 + T25776;
  assign T25776 = $signed(T25777) / $signed(22'h100000);
  assign T25777 = $signed(31'h3da106bd) * $signed(16'h0);
  assign T25778 = {T25781, T25779};
  assign T25779 = $signed(T25780) / $signed(22'h100000);
  assign T25780 = $signed(30'h11423eef) * $signed(16'h1);
  assign T25781 = T25779[6'h2d:6'h2d];
  assign T25782 = T18725[1'h0:1'h0];
  assign T25783 = T18725[1'h1:1'h1];
  assign T25784 = T18725[2'h2:2'h2];
  assign T25785 = T25848 ? T25816 : T25786;
  assign T25786 = T25815 ? T25801 : T25787;
  assign T25787 = T25800 ? twiddle4_1_425_real : twiddle4_1_424_real;
  assign twiddle4_1_424_real = T25790 + T25788;
  assign T25788 = $signed(T25789) / $signed(22'h100000);
  assign T25789 = $signed(31'h3dae81ce) * $signed(16'h0);
  assign T25790 = {T25793, T25791};
  assign T25791 = $signed(T25792) / $signed(22'h100000);
  assign T25792 = $signed(30'h1111d262) * $signed(16'h1);
  assign T25793 = T25791[6'h2d:6'h2d];
  assign twiddle4_1_425_real = T25796 + T25794;
  assign T25794 = $signed(T25795) / $signed(22'h100000);
  assign T25795 = $signed(31'h3dbbd6d4) * $signed(16'h0);
  assign T25796 = {T25799, T25797};
  assign T25797 = $signed(T25798) / $signed(22'h100000);
  assign T25798 = $signed(30'h10e15b4e) * $signed(16'h1);
  assign T25799 = T25797[6'h2d:6'h2d];
  assign T25800 = T18725[1'h0:1'h0];
  assign T25801 = T25814 ? twiddle4_1_427_real : twiddle4_1_426_real;
  assign twiddle4_1_426_real = T25804 + T25802;
  assign T25802 = $signed(T25803) / $signed(22'h100000);
  assign T25803 = $signed(31'h3dc905c4) * $signed(16'h0);
  assign T25804 = {T25807, T25805};
  assign T25805 = $signed(T25806) / $signed(22'h100000);
  assign T25806 = $signed(30'h10b0d9cf) * $signed(16'h1);
  assign T25807 = T25805[6'h2d:6'h2d];
  assign twiddle4_1_427_real = T25810 + T25808;
  assign T25808 = $signed(T25809) / $signed(22'h100000);
  assign T25809 = $signed(31'h3dd60e98) * $signed(16'h0);
  assign T25810 = {T25813, T25811};
  assign T25811 = $signed(T25812) / $signed(22'h100000);
  assign T25812 = $signed(30'h10804e05) * $signed(16'h1);
  assign T25813 = T25811[6'h2d:6'h2d];
  assign T25814 = T18725[1'h0:1'h0];
  assign T25815 = T18725[1'h1:1'h1];
  assign T25816 = T25847 ? T25831 : T25817;
  assign T25817 = T25830 ? twiddle4_1_429_real : twiddle4_1_428_real;
  assign twiddle4_1_428_real = T25820 + T25818;
  assign T25818 = $signed(T25819) / $signed(22'h100000);
  assign T25819 = $signed(31'h3de2f147) * $signed(16'h0);
  assign T25820 = {T25823, T25821};
  assign T25821 = $signed(T25822) / $signed(22'h100000);
  assign T25822 = $signed(30'h104fb80e) * $signed(16'h1);
  assign T25823 = T25821[6'h2d:6'h2d];
  assign twiddle4_1_429_real = T25826 + T25824;
  assign T25824 = $signed(T25825) / $signed(22'h100000);
  assign T25825 = $signed(31'h3defadca) * $signed(16'h0);
  assign T25826 = {T25829, T25827};
  assign T25827 = $signed(T25828) / $signed(22'h100000);
  assign T25828 = $signed(30'h101f1806) * $signed(16'h1);
  assign T25829 = T25827[6'h2d:6'h2d];
  assign T25830 = T18725[1'h0:1'h0];
  assign T25831 = T25846 ? twiddle4_1_431_real : twiddle4_1_430_real;
  assign twiddle4_1_430_real = T25834 + T25832;
  assign T25832 = $signed(T25833) / $signed(22'h100000);
  assign T25833 = $signed(31'h3dfc4418) * $signed(16'h0);
  assign T25834 = {T25837, T25835};
  assign T25835 = $signed(T25836) / $signed(22'h100000);
  assign T25836 = $signed(29'hfee6e0d) * $signed(16'h1);
  assign T25837 = T25838 ? 2'h3 : 2'h0;
  assign T25838 = T25835[6'h2c:6'h2c];
  assign twiddle4_1_431_real = T25841 + T25839;
  assign T25839 = $signed(T25840) / $signed(22'h100000);
  assign T25840 = $signed(31'h3e08b429) * $signed(16'h0);
  assign T25841 = {T25844, T25842};
  assign T25842 = $signed(T25843) / $signed(22'h100000);
  assign T25843 = $signed(29'hfbdba40) * $signed(16'h1);
  assign T25844 = T25845 ? 2'h3 : 2'h0;
  assign T25845 = T25842[6'h2c:6'h2c];
  assign T25846 = T18725[1'h0:1'h0];
  assign T25847 = T18725[1'h1:1'h1];
  assign T25848 = T18725[2'h2:2'h2];
  assign T25849 = T18725[2'h3:2'h3];
  assign T25850 = T25991 ? T25921 : T25851;
  assign T25851 = T25920 ? T25886 : T25852;
  assign T25852 = T25885 ? T25869 : T25853;
  assign T25853 = T25868 ? twiddle4_1_433_real : twiddle4_1_432_real;
  assign twiddle4_1_432_real = T25856 + T25854;
  assign T25854 = $signed(T25855) / $signed(22'h100000);
  assign T25855 = $signed(31'h3e14fdf7) * $signed(16'h0);
  assign T25856 = {T25859, T25857};
  assign T25857 = $signed(T25858) / $signed(22'h100000);
  assign T25858 = $signed(29'hf8cfcbd) * $signed(16'h1);
  assign T25859 = T25860 ? 2'h3 : 2'h0;
  assign T25860 = T25857[6'h2c:6'h2c];
  assign twiddle4_1_433_real = T25863 + T25861;
  assign T25861 = $signed(T25862) / $signed(22'h100000);
  assign T25862 = $signed(31'h3e212179) * $signed(16'h0);
  assign T25863 = {T25866, T25864};
  assign T25864 = $signed(T25865) / $signed(22'h100000);
  assign T25865 = $signed(29'hf5c35a3) * $signed(16'h1);
  assign T25866 = T25867 ? 2'h3 : 2'h0;
  assign T25867 = T25864[6'h2c:6'h2c];
  assign T25868 = T18725[1'h0:1'h0];
  assign T25869 = T25884 ? twiddle4_1_435_real : twiddle4_1_434_real;
  assign twiddle4_1_434_real = T25872 + T25870;
  assign T25870 = $signed(T25871) / $signed(22'h100000);
  assign T25871 = $signed(31'h3e2d1ea7) * $signed(16'h0);
  assign T25872 = {T25875, T25873};
  assign T25873 = $signed(T25874) / $signed(22'h100000);
  assign T25874 = $signed(29'hf2b650f) * $signed(16'h1);
  assign T25875 = T25876 ? 2'h3 : 2'h0;
  assign T25876 = T25873[6'h2c:6'h2c];
  assign twiddle4_1_435_real = T25879 + T25877;
  assign T25877 = $signed(T25878) / $signed(22'h100000);
  assign T25878 = $signed(31'h3e38f57c) * $signed(16'h0);
  assign T25879 = {T25882, T25880};
  assign T25880 = $signed(T25881) / $signed(22'h100000);
  assign T25881 = $signed(29'hefa8b1f) * $signed(16'h1);
  assign T25882 = T25883 ? 2'h3 : 2'h0;
  assign T25883 = T25880[6'h2c:6'h2c];
  assign T25884 = T18725[1'h0:1'h0];
  assign T25885 = T18725[1'h1:1'h1];
  assign T25886 = T25919 ? T25903 : T25887;
  assign T25887 = T25902 ? twiddle4_1_437_real : twiddle4_1_436_real;
  assign twiddle4_1_436_real = T25890 + T25888;
  assign T25888 = $signed(T25889) / $signed(22'h100000);
  assign T25889 = $signed(31'h3e44a5ee) * $signed(16'h0);
  assign T25890 = {T25893, T25891};
  assign T25891 = $signed(T25892) / $signed(22'h100000);
  assign T25892 = $signed(29'hec9a7f2) * $signed(16'h1);
  assign T25893 = T25894 ? 2'h3 : 2'h0;
  assign T25894 = T25891[6'h2c:6'h2c];
  assign twiddle4_1_437_real = T25897 + T25895;
  assign T25895 = $signed(T25896) / $signed(22'h100000);
  assign T25896 = $signed(31'h3e502ff8) * $signed(16'h0);
  assign T25897 = {T25900, T25898};
  assign T25898 = $signed(T25899) / $signed(22'h100000);
  assign T25899 = $signed(29'he98bba6) * $signed(16'h1);
  assign T25900 = T25901 ? 2'h3 : 2'h0;
  assign T25901 = T25898[6'h2c:6'h2c];
  assign T25902 = T18725[1'h0:1'h0];
  assign T25903 = T25918 ? twiddle4_1_439_real : twiddle4_1_438_real;
  assign twiddle4_1_438_real = T25906 + T25904;
  assign T25904 = $signed(T25905) / $signed(22'h100000);
  assign T25905 = $signed(31'h3e5b9392) * $signed(16'h0);
  assign T25906 = {T25909, T25907};
  assign T25907 = $signed(T25908) / $signed(22'h100000);
  assign T25908 = $signed(29'he67c659) * $signed(16'h1);
  assign T25909 = T25910 ? 2'h3 : 2'h0;
  assign T25910 = T25907[6'h2c:6'h2c];
  assign twiddle4_1_439_real = T25913 + T25911;
  assign T25911 = $signed(T25912) / $signed(22'h100000);
  assign T25912 = $signed(31'h3e66d0b4) * $signed(16'h0);
  assign T25913 = {T25916, T25914};
  assign T25914 = $signed(T25915) / $signed(22'h100000);
  assign T25915 = $signed(29'he36c829) * $signed(16'h1);
  assign T25916 = T25917 ? 2'h3 : 2'h0;
  assign T25917 = T25914[6'h2c:6'h2c];
  assign T25918 = T18725[1'h0:1'h0];
  assign T25919 = T18725[1'h1:1'h1];
  assign T25920 = T18725[2'h2:2'h2];
  assign T25921 = T25990 ? T25956 : T25922;
  assign T25922 = T25955 ? T25939 : T25923;
  assign T25923 = T25938 ? twiddle4_1_441_real : twiddle4_1_440_real;
  assign twiddle4_1_440_real = T25926 + T25924;
  assign T25924 = $signed(T25925) / $signed(22'h100000);
  assign T25925 = $signed(31'h3e71e758) * $signed(16'h0);
  assign T25926 = {T25929, T25927};
  assign T25927 = $signed(T25928) / $signed(22'h100000);
  assign T25928 = $signed(29'he05c135) * $signed(16'h1);
  assign T25929 = T25930 ? 2'h3 : 2'h0;
  assign T25930 = T25927[6'h2c:6'h2c];
  assign twiddle4_1_441_real = T25933 + T25931;
  assign T25931 = $signed(T25932) / $signed(22'h100000);
  assign T25932 = $signed(31'h3e7cd778) * $signed(16'h0);
  assign T25933 = {T25936, T25934};
  assign T25934 = $signed(T25935) / $signed(22'h100000);
  assign T25935 = $signed(29'hdd4b19a) * $signed(16'h1);
  assign T25936 = T25937 ? 2'h3 : 2'h0;
  assign T25937 = T25934[6'h2c:6'h2c];
  assign T25938 = T18725[1'h0:1'h0];
  assign T25939 = T25954 ? twiddle4_1_443_real : twiddle4_1_442_real;
  assign twiddle4_1_442_real = T25942 + T25940;
  assign T25940 = $signed(T25941) / $signed(22'h100000);
  assign T25941 = $signed(31'h3e87a10b) * $signed(16'h0);
  assign T25942 = {T25945, T25943};
  assign T25943 = $signed(T25944) / $signed(22'h100000);
  assign T25944 = $signed(29'hda39977) * $signed(16'h1);
  assign T25945 = T25946 ? 2'h3 : 2'h0;
  assign T25946 = T25943[6'h2c:6'h2c];
  assign twiddle4_1_443_real = T25949 + T25947;
  assign T25947 = $signed(T25948) / $signed(22'h100000);
  assign T25948 = $signed(31'h3e92440d) * $signed(16'h0);
  assign T25949 = {T25952, T25950};
  assign T25950 = $signed(T25951) / $signed(22'h100000);
  assign T25951 = $signed(29'hd7278ea) * $signed(16'h1);
  assign T25952 = T25953 ? 2'h3 : 2'h0;
  assign T25953 = T25950[6'h2c:6'h2c];
  assign T25954 = T18725[1'h0:1'h0];
  assign T25955 = T18725[1'h1:1'h1];
  assign T25956 = T25989 ? T25973 : T25957;
  assign T25957 = T25972 ? twiddle4_1_445_real : twiddle4_1_444_real;
  assign twiddle4_1_444_real = T25960 + T25958;
  assign T25958 = $signed(T25959) / $signed(22'h100000);
  assign T25959 = $signed(31'h3e9cc076) * $signed(16'h0);
  assign T25960 = {T25963, T25961};
  assign T25961 = $signed(T25962) / $signed(22'h100000);
  assign T25962 = $signed(29'hd415012) * $signed(16'h1);
  assign T25963 = T25964 ? 2'h3 : 2'h0;
  assign T25964 = T25961[6'h2c:6'h2c];
  assign twiddle4_1_445_real = T25967 + T25965;
  assign T25965 = $signed(T25966) / $signed(22'h100000);
  assign T25966 = $signed(31'h3ea7163f) * $signed(16'h0);
  assign T25967 = {T25970, T25968};
  assign T25968 = $signed(T25969) / $signed(22'h100000);
  assign T25969 = $signed(29'hd101f0d) * $signed(16'h1);
  assign T25970 = T25971 ? 2'h3 : 2'h0;
  assign T25971 = T25968[6'h2c:6'h2c];
  assign T25972 = T18725[1'h0:1'h0];
  assign T25973 = T25988 ? twiddle4_1_447_real : twiddle4_1_446_real;
  assign twiddle4_1_446_real = T25976 + T25974;
  assign T25974 = $signed(T25975) / $signed(22'h100000);
  assign T25975 = $signed(31'h3eb14562) * $signed(16'h0);
  assign T25976 = {T25979, T25977};
  assign T25977 = $signed(T25978) / $signed(22'h100000);
  assign T25978 = $signed(29'hcdee5f9) * $signed(16'h1);
  assign T25979 = T25980 ? 2'h3 : 2'h0;
  assign T25980 = T25977[6'h2c:6'h2c];
  assign twiddle4_1_447_real = T25983 + T25981;
  assign T25981 = $signed(T25982) / $signed(22'h100000);
  assign T25982 = $signed(31'h3ebb4dda) * $signed(16'h0);
  assign T25983 = {T25986, T25984};
  assign T25984 = $signed(T25985) / $signed(22'h100000);
  assign T25985 = $signed(29'hcada4f4) * $signed(16'h1);
  assign T25986 = T25987 ? 2'h3 : 2'h0;
  assign T25987 = T25984[6'h2c:6'h2c];
  assign T25988 = T18725[1'h0:1'h0];
  assign T25989 = T18725[1'h1:1'h1];
  assign T25990 = T18725[2'h2:2'h2];
  assign T25991 = T18725[2'h3:2'h3];
  assign T25992 = T18725[3'h4:3'h4];
  assign T25993 = T18725[3'h5:3'h5];
  assign T25994 = T26567 ? T26281 : T25995;
  assign T25995 = T26280 ? T26138 : T25996;
  assign T25996 = T26137 ? T26067 : T25997;
  assign T25997 = T26066 ? T26032 : T25998;
  assign T25998 = T26031 ? T26015 : T25999;
  assign T25999 = T26014 ? twiddle4_1_449_real : twiddle4_1_448_real;
  assign twiddle4_1_448_real = T26002 + T26000;
  assign T26000 = $signed(T26001) / $signed(22'h100000);
  assign T26001 = $signed(31'h3ec52f9f) * $signed(16'h0);
  assign T26002 = {T26005, T26003};
  assign T26003 = $signed(T26004) / $signed(22'h100000);
  assign T26004 = $signed(29'hc7c5c1e) * $signed(16'h1);
  assign T26005 = T26006 ? 2'h3 : 2'h0;
  assign T26006 = T26003[6'h2c:6'h2c];
  assign twiddle4_1_449_real = T26009 + T26007;
  assign T26007 = $signed(T26008) / $signed(22'h100000);
  assign T26008 = $signed(31'h3eceeaad) * $signed(16'h0);
  assign T26009 = {T26012, T26010};
  assign T26010 = $signed(T26011) / $signed(22'h100000);
  assign T26011 = $signed(29'hc4b0b93) * $signed(16'h1);
  assign T26012 = T26013 ? 2'h3 : 2'h0;
  assign T26013 = T26010[6'h2c:6'h2c];
  assign T26014 = T18725[1'h0:1'h0];
  assign T26015 = T26030 ? twiddle4_1_451_real : twiddle4_1_450_real;
  assign twiddle4_1_450_real = T26018 + T26016;
  assign T26016 = $signed(T26017) / $signed(22'h100000);
  assign T26017 = $signed(31'h3ed87efb) * $signed(16'h0);
  assign T26018 = {T26021, T26019};
  assign T26019 = $signed(T26020) / $signed(22'h100000);
  assign T26020 = $signed(29'hc19b374) * $signed(16'h1);
  assign T26021 = T26022 ? 2'h3 : 2'h0;
  assign T26022 = T26019[6'h2c:6'h2c];
  assign twiddle4_1_451_real = T26025 + T26023;
  assign T26023 = $signed(T26024) / $signed(22'h100000);
  assign T26024 = $signed(31'h3ee1ec86) * $signed(16'h0);
  assign T26025 = {T26028, T26026};
  assign T26026 = $signed(T26027) / $signed(22'h100000);
  assign T26027 = $signed(29'hbe853dd) * $signed(16'h1);
  assign T26028 = T26029 ? 2'h3 : 2'h0;
  assign T26029 = T26026[6'h2c:6'h2c];
  assign T26030 = T18725[1'h0:1'h0];
  assign T26031 = T18725[1'h1:1'h1];
  assign T26032 = T26065 ? T26049 : T26033;
  assign T26033 = T26048 ? twiddle4_1_453_real : twiddle4_1_452_real;
  assign twiddle4_1_452_real = T26036 + T26034;
  assign T26034 = $signed(T26035) / $signed(22'h100000);
  assign T26035 = $signed(31'h3eeb3347) * $signed(16'h0);
  assign T26036 = {T26039, T26037};
  assign T26037 = $signed(T26038) / $signed(22'h100000);
  assign T26038 = $signed(29'hbb6ecef) * $signed(16'h1);
  assign T26039 = T26040 ? 2'h3 : 2'h0;
  assign T26040 = T26037[6'h2c:6'h2c];
  assign twiddle4_1_453_real = T26043 + T26041;
  assign T26041 = $signed(T26042) / $signed(22'h100000);
  assign T26042 = $signed(31'h3ef45338) * $signed(16'h0);
  assign T26043 = {T26046, T26044};
  assign T26044 = $signed(T26045) / $signed(22'h100000);
  assign T26045 = $signed(29'hb857ec6) * $signed(16'h1);
  assign T26046 = T26047 ? 2'h3 : 2'h0;
  assign T26047 = T26044[6'h2c:6'h2c];
  assign T26048 = T18725[1'h0:1'h0];
  assign T26049 = T26064 ? twiddle4_1_455_real : twiddle4_1_454_real;
  assign twiddle4_1_454_real = T26052 + T26050;
  assign T26050 = $signed(T26051) / $signed(22'h100000);
  assign T26051 = $signed(31'h3efd4c53) * $signed(16'h0);
  assign T26052 = {T26055, T26053};
  assign T26053 = $signed(T26054) / $signed(22'h100000);
  assign T26054 = $signed(29'hb540982) * $signed(16'h1);
  assign T26055 = T26056 ? 2'h3 : 2'h0;
  assign T26056 = T26053[6'h2c:6'h2c];
  assign twiddle4_1_455_real = T26059 + T26057;
  assign T26057 = $signed(T26058) / $signed(22'h100000);
  assign T26058 = $signed(31'h3f061e94) * $signed(16'h0);
  assign T26059 = {T26062, T26060};
  assign T26060 = $signed(T26061) / $signed(22'h100000);
  assign T26061 = $signed(29'hb228d41) * $signed(16'h1);
  assign T26062 = T26063 ? 2'h3 : 2'h0;
  assign T26063 = T26060[6'h2c:6'h2c];
  assign T26064 = T18725[1'h0:1'h0];
  assign T26065 = T18725[1'h1:1'h1];
  assign T26066 = T18725[2'h2:2'h2];
  assign T26067 = T26136 ? T26102 : T26068;
  assign T26068 = T26101 ? T26085 : T26069;
  assign T26069 = T26084 ? twiddle4_1_457_real : twiddle4_1_456_real;
  assign twiddle4_1_456_real = T26072 + T26070;
  assign T26070 = $signed(T26071) / $signed(22'h100000);
  assign T26071 = $signed(31'h3f0ec9f4) * $signed(16'h0);
  assign T26072 = {T26075, T26073};
  assign T26073 = $signed(T26074) / $signed(22'h100000);
  assign T26074 = $signed(29'haf10a22) * $signed(16'h1);
  assign T26075 = T26076 ? 2'h3 : 2'h0;
  assign T26076 = T26073[6'h2c:6'h2c];
  assign twiddle4_1_457_real = T26079 + T26077;
  assign T26077 = $signed(T26078) / $signed(22'h100000);
  assign T26078 = $signed(31'h3f174e6f) * $signed(16'h0);
  assign T26079 = {T26082, T26080};
  assign T26080 = $signed(T26081) / $signed(22'h100000);
  assign T26081 = $signed(29'habf8043) * $signed(16'h1);
  assign T26082 = T26083 ? 2'h3 : 2'h0;
  assign T26083 = T26080[6'h2c:6'h2c];
  assign T26084 = T18725[1'h0:1'h0];
  assign T26085 = T26100 ? twiddle4_1_459_real : twiddle4_1_458_real;
  assign twiddle4_1_458_real = T26088 + T26086;
  assign T26086 = $signed(T26087) / $signed(22'h100000);
  assign T26087 = $signed(31'h3f1fabff) * $signed(16'h0);
  assign T26088 = {T26091, T26089};
  assign T26089 = $signed(T26090) / $signed(22'h100000);
  assign T26090 = $signed(29'ha8defc2) * $signed(16'h1);
  assign T26091 = T26092 ? 2'h3 : 2'h0;
  assign T26092 = T26089[6'h2c:6'h2c];
  assign twiddle4_1_459_real = T26095 + T26093;
  assign T26093 = $signed(T26094) / $signed(22'h100000);
  assign T26094 = $signed(31'h3f27e29f) * $signed(16'h0);
  assign T26095 = {T26098, T26096};
  assign T26096 = $signed(T26097) / $signed(22'h100000);
  assign T26097 = $signed(29'ha5c58bf) * $signed(16'h1);
  assign T26098 = T26099 ? 2'h3 : 2'h0;
  assign T26099 = T26096[6'h2c:6'h2c];
  assign T26100 = T18725[1'h0:1'h0];
  assign T26101 = T18725[1'h1:1'h1];
  assign T26102 = T26135 ? T26119 : T26103;
  assign T26103 = T26118 ? twiddle4_1_461_real : twiddle4_1_460_real;
  assign twiddle4_1_460_real = T26106 + T26104;
  assign T26104 = $signed(T26105) / $signed(22'h100000);
  assign T26105 = $signed(31'h3f2ff249) * $signed(16'h0);
  assign T26106 = {T26109, T26107};
  assign T26107 = $signed(T26108) / $signed(22'h100000);
  assign T26108 = $signed(29'ha2abb58) * $signed(16'h1);
  assign T26109 = T26110 ? 2'h3 : 2'h0;
  assign T26110 = T26107[6'h2c:6'h2c];
  assign twiddle4_1_461_real = T26113 + T26111;
  assign T26111 = $signed(T26112) / $signed(22'h100000);
  assign T26112 = $signed(31'h3f37daf9) * $signed(16'h0);
  assign T26113 = {T26116, T26114};
  assign T26114 = $signed(T26115) / $signed(22'h100000);
  assign T26115 = $signed(29'h9f917ab) * $signed(16'h1);
  assign T26116 = T26117 ? 2'h3 : 2'h0;
  assign T26117 = T26114[6'h2c:6'h2c];
  assign T26118 = T18725[1'h0:1'h0];
  assign T26119 = T26134 ? twiddle4_1_463_real : twiddle4_1_462_real;
  assign twiddle4_1_462_real = T26122 + T26120;
  assign T26120 = $signed(T26121) / $signed(22'h100000);
  assign T26121 = $signed(31'h3f3f9cab) * $signed(16'h0);
  assign T26122 = {T26125, T26123};
  assign T26123 = $signed(T26124) / $signed(22'h100000);
  assign T26124 = $signed(29'h9c76dd8) * $signed(16'h1);
  assign T26125 = T26126 ? 2'h3 : 2'h0;
  assign T26126 = T26123[6'h2c:6'h2c];
  assign twiddle4_1_463_real = T26129 + T26127;
  assign T26127 = $signed(T26128) / $signed(22'h100000);
  assign T26128 = $signed(31'h3f473758) * $signed(16'h0);
  assign T26129 = {T26132, T26130};
  assign T26130 = $signed(T26131) / $signed(22'h100000);
  assign T26131 = $signed(29'h995bdfc) * $signed(16'h1);
  assign T26132 = T26133 ? 2'h3 : 2'h0;
  assign T26133 = T26130[6'h2c:6'h2c];
  assign T26134 = T18725[1'h0:1'h0];
  assign T26135 = T18725[1'h1:1'h1];
  assign T26136 = T18725[2'h2:2'h2];
  assign T26137 = T18725[2'h3:2'h3];
  assign T26138 = T26279 ? T26209 : T26139;
  assign T26139 = T26208 ? T26174 : T26140;
  assign T26140 = T26173 ? T26157 : T26141;
  assign T26141 = T26156 ? twiddle4_1_465_real : twiddle4_1_464_real;
  assign twiddle4_1_464_real = T26144 + T26142;
  assign T26142 = $signed(T26143) / $signed(22'h100000);
  assign T26143 = $signed(31'h3f4eaafe) * $signed(16'h0);
  assign T26144 = {T26147, T26145};
  assign T26145 = $signed(T26146) / $signed(22'h100000);
  assign T26146 = $signed(29'h9640837) * $signed(16'h1);
  assign T26147 = T26148 ? 2'h3 : 2'h0;
  assign T26148 = T26145[6'h2c:6'h2c];
  assign twiddle4_1_465_real = T26151 + T26149;
  assign T26149 = $signed(T26150) / $signed(22'h100000);
  assign T26150 = $signed(31'h3f55f796) * $signed(16'h0);
  assign T26151 = {T26154, T26152};
  assign T26152 = $signed(T26153) / $signed(22'h100000);
  assign T26153 = $signed(29'h9324ca6) * $signed(16'h1);
  assign T26154 = T26155 ? 2'h3 : 2'h0;
  assign T26155 = T26152[6'h2c:6'h2c];
  assign T26156 = T18725[1'h0:1'h0];
  assign T26157 = T26172 ? twiddle4_1_467_real : twiddle4_1_466_real;
  assign twiddle4_1_466_real = T26160 + T26158;
  assign T26158 = $signed(T26159) / $signed(22'h100000);
  assign T26159 = $signed(31'h3f5d1d1c) * $signed(16'h0);
  assign T26160 = {T26163, T26161};
  assign T26161 = $signed(T26162) / $signed(22'h100000);
  assign T26162 = $signed(29'h9008b6a) * $signed(16'h1);
  assign T26163 = T26164 ? 2'h3 : 2'h0;
  assign T26164 = T26161[6'h2c:6'h2c];
  assign twiddle4_1_467_real = T26167 + T26165;
  assign T26165 = $signed(T26166) / $signed(22'h100000);
  assign T26166 = $signed(31'h3f641b8d) * $signed(16'h0);
  assign T26167 = {T26170, T26168};
  assign T26168 = $signed(T26169) / $signed(22'h100000);
  assign T26169 = $signed(29'h8cec4a0) * $signed(16'h1);
  assign T26170 = T26171 ? 2'h3 : 2'h0;
  assign T26171 = T26168[6'h2c:6'h2c];
  assign T26172 = T18725[1'h0:1'h0];
  assign T26173 = T18725[1'h1:1'h1];
  assign T26174 = T26207 ? T26191 : T26175;
  assign T26175 = T26190 ? twiddle4_1_469_real : twiddle4_1_468_real;
  assign twiddle4_1_468_real = T26178 + T26176;
  assign T26176 = $signed(T26177) / $signed(22'h100000);
  assign T26177 = $signed(31'h3f6af2e3) * $signed(16'h0);
  assign T26178 = {T26181, T26179};
  assign T26179 = $signed(T26180) / $signed(22'h100000);
  assign T26180 = $signed(29'h89cf867) * $signed(16'h1);
  assign T26181 = T26182 ? 2'h3 : 2'h0;
  assign T26182 = T26179[6'h2c:6'h2c];
  assign twiddle4_1_469_real = T26185 + T26183;
  assign T26183 = $signed(T26184) / $signed(22'h100000);
  assign T26184 = $signed(31'h3f71a31a) * $signed(16'h0);
  assign T26185 = {T26188, T26186};
  assign T26186 = $signed(T26187) / $signed(22'h100000);
  assign T26187 = $signed(29'h86b26de) * $signed(16'h1);
  assign T26188 = T26189 ? 2'h3 : 2'h0;
  assign T26189 = T26186[6'h2c:6'h2c];
  assign T26190 = T18725[1'h0:1'h0];
  assign T26191 = T26206 ? twiddle4_1_471_real : twiddle4_1_470_real;
  assign twiddle4_1_470_real = T26194 + T26192;
  assign T26192 = $signed(T26193) / $signed(22'h100000);
  assign T26193 = $signed(31'h3f782c2f) * $signed(16'h0);
  assign T26194 = {T26197, T26195};
  assign T26195 = $signed(T26196) / $signed(22'h100000);
  assign T26196 = $signed(29'h8395023) * $signed(16'h1);
  assign T26197 = T26198 ? 2'h3 : 2'h0;
  assign T26198 = T26195[6'h2c:6'h2c];
  assign twiddle4_1_471_real = T26201 + T26199;
  assign T26199 = $signed(T26200) / $signed(22'h100000);
  assign T26200 = $signed(31'h3f7e8e1e) * $signed(16'h0);
  assign T26201 = {T26204, T26202};
  assign T26202 = $signed(T26203) / $signed(22'h100000);
  assign T26203 = $signed(29'h8077456) * $signed(16'h1);
  assign T26204 = T26205 ? 2'h3 : 2'h0;
  assign T26205 = T26202[6'h2c:6'h2c];
  assign T26206 = T18725[1'h0:1'h0];
  assign T26207 = T18725[1'h1:1'h1];
  assign T26208 = T18725[2'h2:2'h2];
  assign T26209 = T26278 ? T26244 : T26210;
  assign T26210 = T26243 ? T26227 : T26211;
  assign T26211 = T26226 ? twiddle4_1_473_real : twiddle4_1_472_real;
  assign twiddle4_1_472_real = T26214 + T26212;
  assign T26212 = $signed(T26213) / $signed(22'h100000);
  assign T26213 = $signed(31'h3f84c8e1) * $signed(16'h0);
  assign T26214 = {T26217, T26215};
  assign T26215 = $signed(T26216) / $signed(22'h100000);
  assign T26216 = $signed(28'h7d59395) * $signed(16'h1);
  assign T26217 = T26218 ? 3'h7 : 3'h0;
  assign T26218 = T26215[6'h2b:6'h2b];
  assign twiddle4_1_473_real = T26221 + T26219;
  assign T26219 = $signed(T26220) / $signed(22'h100000);
  assign T26220 = $signed(31'h3f8adc76) * $signed(16'h0);
  assign T26221 = {T26224, T26222};
  assign T26222 = $signed(T26223) / $signed(22'h100000);
  assign T26223 = $signed(28'h7a3adff) * $signed(16'h1);
  assign T26224 = T26225 ? 3'h7 : 3'h0;
  assign T26225 = T26222[6'h2b:6'h2b];
  assign T26226 = T18725[1'h0:1'h0];
  assign T26227 = T26242 ? twiddle4_1_475_real : twiddle4_1_474_real;
  assign twiddle4_1_474_real = T26230 + T26228;
  assign T26228 = $signed(T26229) / $signed(22'h100000);
  assign T26229 = $signed(31'h3f90c8d9) * $signed(16'h0);
  assign T26230 = {T26233, T26231};
  assign T26231 = $signed(T26232) / $signed(22'h100000);
  assign T26232 = $signed(28'h771c3b2) * $signed(16'h1);
  assign T26233 = T26234 ? 3'h7 : 3'h0;
  assign T26234 = T26231[6'h2b:6'h2b];
  assign twiddle4_1_475_real = T26237 + T26235;
  assign T26235 = $signed(T26236) / $signed(22'h100000);
  assign T26236 = $signed(31'h3f968e07) * $signed(16'h0);
  assign T26237 = {T26240, T26238};
  assign T26238 = $signed(T26239) / $signed(22'h100000);
  assign T26239 = $signed(28'h73fd4ce) * $signed(16'h1);
  assign T26240 = T26241 ? 3'h7 : 3'h0;
  assign T26241 = T26238[6'h2b:6'h2b];
  assign T26242 = T18725[1'h0:1'h0];
  assign T26243 = T18725[1'h1:1'h1];
  assign T26244 = T26277 ? T26261 : T26245;
  assign T26245 = T26260 ? twiddle4_1_477_real : twiddle4_1_476_real;
  assign twiddle4_1_476_real = T26248 + T26246;
  assign T26246 = $signed(T26247) / $signed(22'h100000);
  assign T26247 = $signed(31'h3f9c2bfa) * $signed(16'h0);
  assign T26248 = {T26251, T26249};
  assign T26249 = $signed(T26250) / $signed(22'h100000);
  assign T26250 = $signed(28'h70de171) * $signed(16'h1);
  assign T26251 = T26252 ? 3'h7 : 3'h0;
  assign T26252 = T26249[6'h2b:6'h2b];
  assign twiddle4_1_477_real = T26255 + T26253;
  assign T26253 = $signed(T26254) / $signed(22'h100000);
  assign T26254 = $signed(31'h3fa1a2b1) * $signed(16'h0);
  assign T26255 = {T26258, T26256};
  assign T26256 = $signed(T26257) / $signed(22'h100000);
  assign T26257 = $signed(28'h6dbe9bb) * $signed(16'h1);
  assign T26258 = T26259 ? 3'h7 : 3'h0;
  assign T26259 = T26256[6'h2b:6'h2b];
  assign T26260 = T18725[1'h0:1'h0];
  assign T26261 = T26276 ? twiddle4_1_479_real : twiddle4_1_478_real;
  assign twiddle4_1_478_real = T26264 + T26262;
  assign T26262 = $signed(T26263) / $signed(22'h100000);
  assign T26263 = $signed(31'h3fa6f228) * $signed(16'h0);
  assign T26264 = {T26267, T26265};
  assign T26265 = $signed(T26266) / $signed(22'h100000);
  assign T26266 = $signed(28'h6a9edc9) * $signed(16'h1);
  assign T26267 = T26268 ? 3'h7 : 3'h0;
  assign T26268 = T26265[6'h2b:6'h2b];
  assign twiddle4_1_479_real = T26271 + T26269;
  assign T26269 = $signed(T26270) / $signed(22'h100000);
  assign T26270 = $signed(31'h3fac1a5b) * $signed(16'h0);
  assign T26271 = {T26274, T26272};
  assign T26272 = $signed(T26273) / $signed(22'h100000);
  assign T26273 = $signed(28'h677edba) * $signed(16'h1);
  assign T26274 = T26275 ? 3'h7 : 3'h0;
  assign T26275 = T26272[6'h2b:6'h2b];
  assign T26276 = T18725[1'h0:1'h0];
  assign T26277 = T18725[1'h1:1'h1];
  assign T26278 = T18725[2'h2:2'h2];
  assign T26279 = T18725[2'h3:2'h3];
  assign T26280 = T18725[3'h4:3'h4];
  assign T26281 = T26566 ? T26424 : T26282;
  assign T26282 = T26423 ? T26353 : T26283;
  assign T26283 = T26352 ? T26318 : T26284;
  assign T26284 = T26317 ? T26301 : T26285;
  assign T26285 = T26300 ? twiddle4_1_481_real : twiddle4_1_480_real;
  assign twiddle4_1_480_real = T26288 + T26286;
  assign T26286 = $signed(T26287) / $signed(22'h100000);
  assign T26287 = $signed(31'h3fb11b47) * $signed(16'h0);
  assign T26288 = {T26291, T26289};
  assign T26289 = $signed(T26290) / $signed(22'h100000);
  assign T26290 = $signed(28'h645e9af) * $signed(16'h1);
  assign T26291 = T26292 ? 3'h7 : 3'h0;
  assign T26292 = T26289[6'h2b:6'h2b];
  assign twiddle4_1_481_real = T26295 + T26293;
  assign T26293 = $signed(T26294) / $signed(22'h100000);
  assign T26294 = $signed(31'h3fb5f4ea) * $signed(16'h0);
  assign T26295 = {T26298, T26296};
  assign T26296 = $signed(T26297) / $signed(22'h100000);
  assign T26297 = $signed(28'h613e1c4) * $signed(16'h1);
  assign T26298 = T26299 ? 3'h7 : 3'h0;
  assign T26299 = T26296[6'h2b:6'h2b];
  assign T26300 = T18725[1'h0:1'h0];
  assign T26301 = T26316 ? twiddle4_1_483_real : twiddle4_1_482_real;
  assign twiddle4_1_482_real = T26304 + T26302;
  assign T26302 = $signed(T26303) / $signed(22'h100000);
  assign T26303 = $signed(31'h3fbaa73f) * $signed(16'h0);
  assign T26304 = {T26307, T26305};
  assign T26305 = $signed(T26306) / $signed(22'h100000);
  assign T26306 = $signed(28'h5e1d61a) * $signed(16'h1);
  assign T26307 = T26308 ? 3'h7 : 3'h0;
  assign T26308 = T26305[6'h2b:6'h2b];
  assign twiddle4_1_483_real = T26311 + T26309;
  assign T26309 = $signed(T26310) / $signed(22'h100000);
  assign T26310 = $signed(31'h3fbf3245) * $signed(16'h0);
  assign T26311 = {T26314, T26312};
  assign T26312 = $signed(T26313) / $signed(22'h100000);
  assign T26313 = $signed(28'h5afc6cf) * $signed(16'h1);
  assign T26314 = T26315 ? 3'h7 : 3'h0;
  assign T26315 = T26312[6'h2b:6'h2b];
  assign T26316 = T18725[1'h0:1'h0];
  assign T26317 = T18725[1'h1:1'h1];
  assign T26318 = T26351 ? T26335 : T26319;
  assign T26319 = T26334 ? twiddle4_1_485_real : twiddle4_1_484_real;
  assign twiddle4_1_484_real = T26322 + T26320;
  assign T26320 = $signed(T26321) / $signed(22'h100000);
  assign T26321 = $signed(31'h3fc395f9) * $signed(16'h0);
  assign T26322 = {T26325, T26323};
  assign T26323 = $signed(T26324) / $signed(22'h100000);
  assign T26324 = $signed(28'h57db402) * $signed(16'h1);
  assign T26325 = T26326 ? 3'h7 : 3'h0;
  assign T26326 = T26323[6'h2b:6'h2b];
  assign twiddle4_1_485_real = T26329 + T26327;
  assign T26327 = $signed(T26328) / $signed(22'h100000);
  assign T26328 = $signed(31'h3fc7d257) * $signed(16'h0);
  assign T26329 = {T26332, T26330};
  assign T26330 = $signed(T26331) / $signed(22'h100000);
  assign T26331 = $signed(28'h54b9dd2) * $signed(16'h1);
  assign T26332 = T26333 ? 3'h7 : 3'h0;
  assign T26333 = T26330[6'h2b:6'h2b];
  assign T26334 = T18725[1'h0:1'h0];
  assign T26335 = T26350 ? twiddle4_1_487_real : twiddle4_1_486_real;
  assign twiddle4_1_486_real = T26338 + T26336;
  assign T26336 = $signed(T26337) / $signed(22'h100000);
  assign T26337 = $signed(31'h3fcbe75e) * $signed(16'h0);
  assign T26338 = {T26341, T26339};
  assign T26339 = $signed(T26340) / $signed(22'h100000);
  assign T26340 = $signed(28'h519845e) * $signed(16'h1);
  assign T26341 = T26342 ? 3'h7 : 3'h0;
  assign T26342 = T26339[6'h2b:6'h2b];
  assign twiddle4_1_487_real = T26345 + T26343;
  assign T26343 = $signed(T26344) / $signed(22'h100000);
  assign T26344 = $signed(31'h3fcfd50a) * $signed(16'h0);
  assign T26345 = {T26348, T26346};
  assign T26346 = $signed(T26347) / $signed(22'h100000);
  assign T26347 = $signed(28'h4e767c4) * $signed(16'h1);
  assign T26348 = T26349 ? 3'h7 : 3'h0;
  assign T26349 = T26346[6'h2b:6'h2b];
  assign T26350 = T18725[1'h0:1'h0];
  assign T26351 = T18725[1'h1:1'h1];
  assign T26352 = T18725[2'h2:2'h2];
  assign T26353 = T26422 ? T26388 : T26354;
  assign T26354 = T26387 ? T26371 : T26355;
  assign T26355 = T26370 ? twiddle4_1_489_real : twiddle4_1_488_real;
  assign twiddle4_1_488_real = T26358 + T26356;
  assign T26356 = $signed(T26357) / $signed(22'h100000);
  assign T26357 = $signed(31'h3fd39b5a) * $signed(16'h0);
  assign T26358 = {T26361, T26359};
  assign T26359 = $signed(T26360) / $signed(22'h100000);
  assign T26360 = $signed(28'h4b54824) * $signed(16'h1);
  assign T26361 = T26362 ? 3'h7 : 3'h0;
  assign T26362 = T26359[6'h2b:6'h2b];
  assign twiddle4_1_489_real = T26365 + T26363;
  assign T26363 = $signed(T26364) / $signed(22'h100000);
  assign T26364 = $signed(31'h3fd73a4a) * $signed(16'h0);
  assign T26365 = {T26368, T26366};
  assign T26366 = $signed(T26367) / $signed(22'h100000);
  assign T26367 = $signed(28'h483259d) * $signed(16'h1);
  assign T26368 = T26369 ? 3'h7 : 3'h0;
  assign T26369 = T26366[6'h2b:6'h2b];
  assign T26370 = T18725[1'h0:1'h0];
  assign T26371 = T26386 ? twiddle4_1_491_real : twiddle4_1_490_real;
  assign twiddle4_1_490_real = T26374 + T26372;
  assign T26372 = $signed(T26373) / $signed(22'h100000);
  assign T26373 = $signed(31'h3fdab1d9) * $signed(16'h0);
  assign T26374 = {T26377, T26375};
  assign T26375 = $signed(T26376) / $signed(22'h100000);
  assign T26376 = $signed(28'h451004d) * $signed(16'h1);
  assign T26377 = T26378 ? 3'h7 : 3'h0;
  assign T26378 = T26375[6'h2b:6'h2b];
  assign twiddle4_1_491_real = T26381 + T26379;
  assign T26379 = $signed(T26380) / $signed(22'h100000);
  assign T26380 = $signed(31'h3fde0205) * $signed(16'h0);
  assign T26381 = {T26384, T26382};
  assign T26382 = $signed(T26383) / $signed(22'h100000);
  assign T26383 = $signed(28'h41ed853) * $signed(16'h1);
  assign T26384 = T26385 ? 3'h7 : 3'h0;
  assign T26385 = T26382[6'h2b:6'h2b];
  assign T26386 = T18725[1'h0:1'h0];
  assign T26387 = T18725[1'h1:1'h1];
  assign T26388 = T26421 ? T26405 : T26389;
  assign T26389 = T26404 ? twiddle4_1_493_real : twiddle4_1_492_real;
  assign twiddle4_1_492_real = T26392 + T26390;
  assign T26390 = $signed(T26391) / $signed(22'h100000);
  assign T26391 = $signed(31'h3fe12acb) * $signed(16'h0);
  assign T26392 = {T26395, T26393};
  assign T26393 = $signed(T26394) / $signed(22'h100000);
  assign T26394 = $signed(27'h3ecadcf) * $signed(16'h1);
  assign T26395 = T26396 ? 4'hf : 4'h0;
  assign T26396 = T26393[6'h2a:6'h2a];
  assign twiddle4_1_493_real = T26399 + T26397;
  assign T26397 = $signed(T26398) / $signed(22'h100000);
  assign T26398 = $signed(31'h3fe42c29) * $signed(16'h0);
  assign T26399 = {T26402, T26400};
  assign T26400 = $signed(T26401) / $signed(22'h100000);
  assign T26401 = $signed(27'h3ba80df) * $signed(16'h1);
  assign T26402 = T26403 ? 4'hf : 4'h0;
  assign T26403 = T26400[6'h2a:6'h2a];
  assign T26404 = T18725[1'h0:1'h0];
  assign T26405 = T26420 ? twiddle4_1_495_real : twiddle4_1_494_real;
  assign twiddle4_1_494_real = T26408 + T26406;
  assign T26406 = $signed(T26407) / $signed(22'h100000);
  assign T26407 = $signed(31'h3fe7061f) * $signed(16'h0);
  assign T26408 = {T26411, T26409};
  assign T26409 = $signed(T26410) / $signed(22'h100000);
  assign T26410 = $signed(27'h38851a2) * $signed(16'h1);
  assign T26411 = T26412 ? 4'hf : 4'h0;
  assign T26412 = T26409[6'h2a:6'h2a];
  assign twiddle4_1_495_real = T26415 + T26413;
  assign T26413 = $signed(T26414) / $signed(22'h100000);
  assign T26414 = $signed(31'h3fe9b8a9) * $signed(16'h0);
  assign T26415 = {T26418, T26416};
  assign T26416 = $signed(T26417) / $signed(22'h100000);
  assign T26417 = $signed(27'h3562037) * $signed(16'h1);
  assign T26418 = T26419 ? 4'hf : 4'h0;
  assign T26419 = T26416[6'h2a:6'h2a];
  assign T26420 = T18725[1'h0:1'h0];
  assign T26421 = T18725[1'h1:1'h1];
  assign T26422 = T18725[2'h2:2'h2];
  assign T26423 = T18725[2'h3:2'h3];
  assign T26424 = T26565 ? T26495 : T26425;
  assign T26425 = T26494 ? T26460 : T26426;
  assign T26426 = T26459 ? T26443 : T26427;
  assign T26427 = T26442 ? twiddle4_1_497_real : twiddle4_1_496_real;
  assign twiddle4_1_496_real = T26430 + T26428;
  assign T26428 = $signed(T26429) / $signed(22'h100000);
  assign T26429 = $signed(31'h3fec43c6) * $signed(16'h0);
  assign T26430 = {T26433, T26431};
  assign T26431 = $signed(T26432) / $signed(22'h100000);
  assign T26432 = $signed(27'h323ecbe) * $signed(16'h1);
  assign T26433 = T26434 ? 4'hf : 4'h0;
  assign T26434 = T26431[6'h2a:6'h2a];
  assign twiddle4_1_497_real = T26437 + T26435;
  assign T26435 = $signed(T26436) / $signed(22'h100000);
  assign T26436 = $signed(31'h3feea776) * $signed(16'h0);
  assign T26437 = {T26440, T26438};
  assign T26438 = $signed(T26439) / $signed(22'h100000);
  assign T26439 = $signed(27'h2f1b754) * $signed(16'h1);
  assign T26440 = T26441 ? 4'hf : 4'h0;
  assign T26441 = T26438[6'h2a:6'h2a];
  assign T26442 = T18725[1'h0:1'h0];
  assign T26443 = T26458 ? twiddle4_1_499_real : twiddle4_1_498_real;
  assign twiddle4_1_498_real = T26446 + T26444;
  assign T26444 = $signed(T26445) / $signed(22'h100000);
  assign T26445 = $signed(31'h3ff0e3b5) * $signed(16'h0);
  assign T26446 = {T26449, T26447};
  assign T26447 = $signed(T26448) / $signed(22'h100000);
  assign T26448 = $signed(27'h2bf801a) * $signed(16'h1);
  assign T26449 = T26450 ? 4'hf : 4'h0;
  assign T26450 = T26447[6'h2a:6'h2a];
  assign twiddle4_1_499_real = T26453 + T26451;
  assign T26451 = $signed(T26452) / $signed(22'h100000);
  assign T26452 = $signed(31'h3ff2f884) * $signed(16'h0);
  assign T26453 = {T26456, T26454};
  assign T26454 = $signed(T26455) / $signed(22'h100000);
  assign T26455 = $signed(27'h28d472d) * $signed(16'h1);
  assign T26456 = T26457 ? 4'hf : 4'h0;
  assign T26457 = T26454[6'h2a:6'h2a];
  assign T26458 = T18725[1'h0:1'h0];
  assign T26459 = T18725[1'h1:1'h1];
  assign T26460 = T26493 ? T26477 : T26461;
  assign T26461 = T26476 ? twiddle4_1_501_real : twiddle4_1_500_real;
  assign twiddle4_1_500_real = T26464 + T26462;
  assign T26462 = $signed(T26463) / $signed(22'h100000);
  assign T26463 = $signed(31'h3ff4e5df) * $signed(16'h0);
  assign T26464 = {T26467, T26465};
  assign T26465 = $signed(T26466) / $signed(22'h100000);
  assign T26466 = $signed(27'h25b0cae) * $signed(16'h1);
  assign T26467 = T26468 ? 4'hf : 4'h0;
  assign T26468 = T26465[6'h2a:6'h2a];
  assign twiddle4_1_501_real = T26471 + T26469;
  assign T26469 = $signed(T26470) / $signed(22'h100000);
  assign T26470 = $signed(31'h3ff6abc8) * $signed(16'h0);
  assign T26471 = {T26474, T26472};
  assign T26472 = $signed(T26473) / $signed(22'h100000);
  assign T26473 = $signed(27'h228d0bb) * $signed(16'h1);
  assign T26474 = T26475 ? 4'hf : 4'h0;
  assign T26475 = T26472[6'h2a:6'h2a];
  assign T26476 = T18725[1'h0:1'h0];
  assign T26477 = T26492 ? twiddle4_1_503_real : twiddle4_1_502_real;
  assign twiddle4_1_502_real = T26480 + T26478;
  assign T26478 = $signed(T26479) / $signed(22'h100000);
  assign T26479 = $signed(31'h3ff84a3b) * $signed(16'h0);
  assign T26480 = {T26483, T26481};
  assign T26481 = $signed(T26482) / $signed(22'h100000);
  assign T26482 = $signed(26'h1f69373) * $signed(16'h1);
  assign T26483 = T26484 ? 5'h1f : 5'h0;
  assign T26484 = T26481[6'h29:6'h29];
  assign twiddle4_1_503_real = T26487 + T26485;
  assign T26485 = $signed(T26486) / $signed(22'h100000);
  assign T26486 = $signed(31'h3ff9c139) * $signed(16'h0);
  assign T26487 = {T26490, T26488};
  assign T26488 = $signed(T26489) / $signed(22'h100000);
  assign T26489 = $signed(26'h1c454f4) * $signed(16'h1);
  assign T26490 = T26491 ? 5'h1f : 5'h0;
  assign T26491 = T26488[6'h29:6'h29];
  assign T26492 = T18725[1'h0:1'h0];
  assign T26493 = T18725[1'h1:1'h1];
  assign T26494 = T18725[2'h2:2'h2];
  assign T26495 = T26564 ? T26530 : T26496;
  assign T26496 = T26529 ? T26513 : T26497;
  assign T26497 = T26512 ? twiddle4_1_505_real : twiddle4_1_504_real;
  assign twiddle4_1_504_real = T26500 + T26498;
  assign T26498 = $signed(T26499) / $signed(22'h100000);
  assign T26499 = $signed(31'h3ffb10c1) * $signed(16'h0);
  assign T26500 = {T26503, T26501};
  assign T26501 = $signed(T26502) / $signed(22'h100000);
  assign T26502 = $signed(26'h192155f) * $signed(16'h1);
  assign T26503 = T26504 ? 5'h1f : 5'h0;
  assign T26504 = T26501[6'h29:6'h29];
  assign twiddle4_1_505_real = T26507 + T26505;
  assign T26505 = $signed(T26506) / $signed(22'h100000);
  assign T26506 = $signed(31'h3ffc38d0) * $signed(16'h0);
  assign T26507 = {T26510, T26508};
  assign T26508 = $signed(T26509) / $signed(22'h100000);
  assign T26509 = $signed(26'h15fd4d2) * $signed(16'h1);
  assign T26510 = T26511 ? 5'h1f : 5'h0;
  assign T26511 = T26508[6'h29:6'h29];
  assign T26512 = T18725[1'h0:1'h0];
  assign T26513 = T26528 ? twiddle4_1_507_real : twiddle4_1_506_real;
  assign twiddle4_1_506_real = T26516 + T26514;
  assign T26514 = $signed(T26515) / $signed(22'h100000);
  assign T26515 = $signed(31'h3ffd3968) * $signed(16'h0);
  assign T26516 = {T26519, T26517};
  assign T26517 = $signed(T26518) / $signed(22'h100000);
  assign T26518 = $signed(26'h12d936b) * $signed(16'h1);
  assign T26519 = T26520 ? 5'h1f : 5'h0;
  assign T26520 = T26517[6'h29:6'h29];
  assign twiddle4_1_507_real = T26523 + T26521;
  assign T26521 = $signed(T26522) / $signed(22'h100000);
  assign T26522 = $signed(31'h3ffe1287) * $signed(16'h0);
  assign T26523 = {T26526, T26524};
  assign T26524 = $signed(T26525) / $signed(22'h100000);
  assign T26525 = $signed(25'hfb514b) * $signed(16'h1);
  assign T26526 = T26527 ? 6'h3f : 6'h0;
  assign T26527 = T26524[6'h28:6'h28];
  assign T26528 = T18725[1'h0:1'h0];
  assign T26529 = T18725[1'h1:1'h1];
  assign T26530 = T26563 ? T26547 : T26531;
  assign T26531 = T26546 ? twiddle4_1_509_real : twiddle4_1_508_real;
  assign twiddle4_1_508_real = T26534 + T26532;
  assign T26532 = $signed(T26533) / $signed(22'h100000);
  assign T26533 = $signed(31'h3ffec42d) * $signed(16'h0);
  assign T26534 = {T26537, T26535};
  assign T26535 = $signed(T26536) / $signed(22'h100000);
  assign T26536 = $signed(25'hc90e8f) * $signed(16'h1);
  assign T26537 = T26538 ? 6'h3f : 6'h0;
  assign T26538 = T26535[6'h28:6'h28];
  assign twiddle4_1_509_real = T26541 + T26539;
  assign T26539 = $signed(T26540) / $signed(22'h100000);
  assign T26540 = $signed(31'h3fff4e59) * $signed(16'h0);
  assign T26541 = {T26544, T26542};
  assign T26542 = $signed(T26543) / $signed(22'h100000);
  assign T26543 = $signed(25'h96cb58) * $signed(16'h1);
  assign T26544 = T26545 ? 6'h3f : 6'h0;
  assign T26545 = T26542[6'h28:6'h28];
  assign T26546 = T18725[1'h0:1'h0];
  assign T26547 = T26562 ? twiddle4_1_511_real : twiddle4_1_510_real;
  assign twiddle4_1_510_real = T26550 + T26548;
  assign T26548 = $signed(T26549) / $signed(22'h100000);
  assign T26549 = $signed(31'h3fffb10b) * $signed(16'h0);
  assign T26550 = {T26553, T26551};
  assign T26551 = $signed(T26552) / $signed(22'h100000);
  assign T26552 = $signed(24'h6487c3) * $signed(16'h1);
  assign T26553 = T26554 ? 7'h7f : 7'h0;
  assign T26554 = T26551[6'h27:6'h27];
  assign twiddle4_1_511_real = T26557 + T26555;
  assign T26555 = $signed(T26556) / $signed(22'h100000);
  assign T26556 = $signed(31'h3fffec42) * $signed(16'h0);
  assign T26557 = {T26560, T26558};
  assign T26558 = $signed(T26559) / $signed(22'h100000);
  assign T26559 = $signed(23'h3243f1) * $signed(16'h1);
  assign T26560 = T26561 ? 8'hff : 8'h0;
  assign T26561 = T26558[6'h26:6'h26];
  assign T26562 = T18725[1'h0:1'h0];
  assign T26563 = T18725[1'h1:1'h1];
  assign T26564 = T18725[2'h2:2'h2];
  assign T26565 = T18725[2'h3:2'h3];
  assign T26566 = T18725[3'h4:3'h4];
  assign T26567 = T18725[3'h5:3'h5];
  assign T26568 = T18725[3'h6:3'h6];
  assign T26569 = T18725[3'h7:3'h7];
  assign T26570 = T24614[6'h2e:6'h2e];
  assign T26571 = T18725[4'h8:4'h8];
endmodule

