module r3icLUT(
    input [10:0] io_ina,
    input [2:0] io_inb,
    output[2:0] io_r3IC
);

  wire[2:0] T0;
  wire[1:0] T1;
  reg [1:0] T2 [1214:0];
  wire[10:0] T3;
  wire[13:0] T4;
  wire[13:0] T5;
  wire[13:0] index;


  assign io_r3IC = T0;
  assign T0 = {1'h0, T1};
`ifndef SYNTHESIS
  assign T1 = T3 >= 11'h4bf ? {1{$random}} : T2[T3];
`else
  assign T1 = T2[T3];
`endif
  always @(*) begin
    T2[0] = 2'h0;
    T2[1] = 2'h0;
    T2[2] = 2'h0;
    T2[3] = 2'h0;
    T2[4] = 2'h0;
    T2[5] = 2'h1;
    T2[6] = 2'h0;
    T2[7] = 2'h0;
    T2[8] = 2'h0;
    T2[9] = 2'h0;
    T2[10] = 2'h2;
    T2[11] = 2'h0;
    T2[12] = 2'h0;
    T2[13] = 2'h0;
    T2[14] = 2'h0;
    T2[15] = 2'h0;
    T2[16] = 2'h1;
    T2[17] = 2'h0;
    T2[18] = 2'h0;
    T2[19] = 2'h0;
    T2[20] = 2'h1;
    T2[21] = 2'h1;
    T2[22] = 2'h0;
    T2[23] = 2'h0;
    T2[24] = 2'h0;
    T2[25] = 2'h2;
    T2[26] = 2'h1;
    T2[27] = 2'h0;
    T2[28] = 2'h0;
    T2[29] = 2'h0;
    T2[30] = 2'h0;
    T2[31] = 2'h2;
    T2[32] = 2'h0;
    T2[33] = 2'h0;
    T2[34] = 2'h0;
    T2[35] = 2'h1;
    T2[36] = 2'h2;
    T2[37] = 2'h0;
    T2[38] = 2'h0;
    T2[39] = 2'h0;
    T2[40] = 2'h2;
    T2[41] = 2'h2;
    T2[42] = 2'h0;
    T2[43] = 2'h0;
    T2[44] = 2'h0;
    T2[45] = 2'h0;
    T2[46] = 2'h0;
    T2[47] = 2'h1;
    T2[48] = 2'h0;
    T2[49] = 2'h0;
    T2[50] = 2'h1;
    T2[51] = 2'h0;
    T2[52] = 2'h1;
    T2[53] = 2'h0;
    T2[54] = 2'h0;
    T2[55] = 2'h2;
    T2[56] = 2'h0;
    T2[57] = 2'h1;
    T2[58] = 2'h0;
    T2[59] = 2'h0;
    T2[60] = 2'h0;
    T2[61] = 2'h1;
    T2[62] = 2'h1;
    T2[63] = 2'h0;
    T2[64] = 2'h0;
    T2[65] = 2'h1;
    T2[66] = 2'h1;
    T2[67] = 2'h1;
    T2[68] = 2'h0;
    T2[69] = 2'h0;
    T2[70] = 2'h2;
    T2[71] = 2'h1;
    T2[72] = 2'h1;
    T2[73] = 2'h0;
    T2[74] = 2'h0;
    T2[75] = 2'h0;
    T2[76] = 2'h2;
    T2[77] = 2'h1;
    T2[78] = 2'h0;
    T2[79] = 2'h0;
    T2[80] = 2'h1;
    T2[81] = 2'h2;
    T2[82] = 2'h1;
    T2[83] = 2'h0;
    T2[84] = 2'h0;
    T2[85] = 2'h2;
    T2[86] = 2'h2;
    T2[87] = 2'h1;
    T2[88] = 2'h0;
    T2[89] = 2'h0;
    T2[90] = 2'h0;
    T2[91] = 2'h0;
    T2[92] = 2'h2;
    T2[93] = 2'h0;
    T2[94] = 2'h0;
    T2[95] = 2'h1;
    T2[96] = 2'h0;
    T2[97] = 2'h2;
    T2[98] = 2'h0;
    T2[99] = 2'h0;
    T2[100] = 2'h2;
    T2[101] = 2'h0;
    T2[102] = 2'h2;
    T2[103] = 2'h0;
    T2[104] = 2'h0;
    T2[105] = 2'h0;
    T2[106] = 2'h1;
    T2[107] = 2'h2;
    T2[108] = 2'h0;
    T2[109] = 2'h0;
    T2[110] = 2'h1;
    T2[111] = 2'h1;
    T2[112] = 2'h2;
    T2[113] = 2'h0;
    T2[114] = 2'h0;
    T2[115] = 2'h2;
    T2[116] = 2'h1;
    T2[117] = 2'h2;
    T2[118] = 2'h0;
    T2[119] = 2'h0;
    T2[120] = 2'h0;
    T2[121] = 2'h2;
    T2[122] = 2'h2;
    T2[123] = 2'h0;
    T2[124] = 2'h0;
    T2[125] = 2'h1;
    T2[126] = 2'h2;
    T2[127] = 2'h2;
    T2[128] = 2'h0;
    T2[129] = 2'h0;
    T2[130] = 2'h2;
    T2[131] = 2'h2;
    T2[132] = 2'h2;
    T2[133] = 2'h0;
    T2[134] = 2'h0;
    T2[135] = 2'h0;
    T2[136] = 2'h0;
    T2[137] = 2'h0;
    T2[138] = 2'h1;
    T2[139] = 2'h0;
    T2[140] = 2'h1;
    T2[141] = 2'h0;
    T2[142] = 2'h0;
    T2[143] = 2'h1;
    T2[144] = 2'h0;
    T2[145] = 2'h2;
    T2[146] = 2'h0;
    T2[147] = 2'h0;
    T2[148] = 2'h1;
    T2[149] = 2'h0;
    T2[150] = 2'h0;
    T2[151] = 2'h1;
    T2[152] = 2'h0;
    T2[153] = 2'h1;
    T2[154] = 2'h0;
    T2[155] = 2'h1;
    T2[156] = 2'h1;
    T2[157] = 2'h0;
    T2[158] = 2'h1;
    T2[159] = 2'h0;
    T2[160] = 2'h2;
    T2[161] = 2'h1;
    T2[162] = 2'h0;
    T2[163] = 2'h1;
    T2[164] = 2'h0;
    T2[165] = 2'h0;
    T2[166] = 2'h2;
    T2[167] = 2'h0;
    T2[168] = 2'h1;
    T2[169] = 2'h0;
    T2[170] = 2'h1;
    T2[171] = 2'h2;
    T2[172] = 2'h0;
    T2[173] = 2'h1;
    T2[174] = 2'h0;
    T2[175] = 2'h2;
    T2[176] = 2'h2;
    T2[177] = 2'h0;
    T2[178] = 2'h1;
    T2[179] = 2'h0;
    T2[180] = 2'h0;
    T2[181] = 2'h0;
    T2[182] = 2'h1;
    T2[183] = 2'h1;
    T2[184] = 2'h0;
    T2[185] = 2'h1;
    T2[186] = 2'h0;
    T2[187] = 2'h1;
    T2[188] = 2'h1;
    T2[189] = 2'h0;
    T2[190] = 2'h2;
    T2[191] = 2'h0;
    T2[192] = 2'h1;
    T2[193] = 2'h1;
    T2[194] = 2'h0;
    T2[195] = 2'h0;
    T2[196] = 2'h1;
    T2[197] = 2'h1;
    T2[198] = 2'h1;
    T2[199] = 2'h0;
    T2[200] = 2'h1;
    T2[201] = 2'h1;
    T2[202] = 2'h1;
    T2[203] = 2'h1;
    T2[204] = 2'h0;
    T2[205] = 2'h2;
    T2[206] = 2'h1;
    T2[207] = 2'h1;
    T2[208] = 2'h1;
    T2[209] = 2'h0;
    T2[210] = 2'h0;
    T2[211] = 2'h2;
    T2[212] = 2'h1;
    T2[213] = 2'h1;
    T2[214] = 2'h0;
    T2[215] = 2'h1;
    T2[216] = 2'h2;
    T2[217] = 2'h1;
    T2[218] = 2'h1;
    T2[219] = 2'h0;
    T2[220] = 2'h2;
    T2[221] = 2'h2;
    T2[222] = 2'h1;
    T2[223] = 2'h1;
    T2[224] = 2'h0;
    T2[225] = 2'h0;
    T2[226] = 2'h0;
    T2[227] = 2'h2;
    T2[228] = 2'h1;
    T2[229] = 2'h0;
    T2[230] = 2'h1;
    T2[231] = 2'h0;
    T2[232] = 2'h2;
    T2[233] = 2'h1;
    T2[234] = 2'h0;
    T2[235] = 2'h2;
    T2[236] = 2'h0;
    T2[237] = 2'h2;
    T2[238] = 2'h1;
    T2[239] = 2'h0;
    T2[240] = 2'h0;
    T2[241] = 2'h1;
    T2[242] = 2'h2;
    T2[243] = 2'h1;
    T2[244] = 2'h0;
    T2[245] = 2'h1;
    T2[246] = 2'h1;
    T2[247] = 2'h2;
    T2[248] = 2'h1;
    T2[249] = 2'h0;
    T2[250] = 2'h2;
    T2[251] = 2'h1;
    T2[252] = 2'h2;
    T2[253] = 2'h1;
    T2[254] = 2'h0;
    T2[255] = 2'h0;
    T2[256] = 2'h2;
    T2[257] = 2'h2;
    T2[258] = 2'h1;
    T2[259] = 2'h0;
    T2[260] = 2'h1;
    T2[261] = 2'h2;
    T2[262] = 2'h2;
    T2[263] = 2'h1;
    T2[264] = 2'h0;
    T2[265] = 2'h2;
    T2[266] = 2'h2;
    T2[267] = 2'h2;
    T2[268] = 2'h1;
    T2[269] = 2'h0;
    T2[270] = 2'h0;
    T2[271] = 2'h0;
    T2[272] = 2'h0;
    T2[273] = 2'h2;
    T2[274] = 2'h0;
    T2[275] = 2'h1;
    T2[276] = 2'h0;
    T2[277] = 2'h0;
    T2[278] = 2'h2;
    T2[279] = 2'h0;
    T2[280] = 2'h2;
    T2[281] = 2'h0;
    T2[282] = 2'h0;
    T2[283] = 2'h2;
    T2[284] = 2'h0;
    T2[285] = 2'h0;
    T2[286] = 2'h1;
    T2[287] = 2'h0;
    T2[288] = 2'h2;
    T2[289] = 2'h0;
    T2[290] = 2'h1;
    T2[291] = 2'h1;
    T2[292] = 2'h0;
    T2[293] = 2'h2;
    T2[294] = 2'h0;
    T2[295] = 2'h2;
    T2[296] = 2'h1;
    T2[297] = 2'h0;
    T2[298] = 2'h2;
    T2[299] = 2'h0;
    T2[300] = 2'h0;
    T2[301] = 2'h2;
    T2[302] = 2'h0;
    T2[303] = 2'h2;
    T2[304] = 2'h0;
    T2[305] = 2'h1;
    T2[306] = 2'h2;
    T2[307] = 2'h0;
    T2[308] = 2'h2;
    T2[309] = 2'h0;
    T2[310] = 2'h2;
    T2[311] = 2'h2;
    T2[312] = 2'h0;
    T2[313] = 2'h2;
    T2[314] = 2'h0;
    T2[315] = 2'h0;
    T2[316] = 2'h0;
    T2[317] = 2'h1;
    T2[318] = 2'h2;
    T2[319] = 2'h0;
    T2[320] = 2'h1;
    T2[321] = 2'h0;
    T2[322] = 2'h1;
    T2[323] = 2'h2;
    T2[324] = 2'h0;
    T2[325] = 2'h2;
    T2[326] = 2'h0;
    T2[327] = 2'h1;
    T2[328] = 2'h2;
    T2[329] = 2'h0;
    T2[330] = 2'h0;
    T2[331] = 2'h1;
    T2[332] = 2'h1;
    T2[333] = 2'h2;
    T2[334] = 2'h0;
    T2[335] = 2'h1;
    T2[336] = 2'h1;
    T2[337] = 2'h1;
    T2[338] = 2'h2;
    T2[339] = 2'h0;
    T2[340] = 2'h2;
    T2[341] = 2'h1;
    T2[342] = 2'h1;
    T2[343] = 2'h2;
    T2[344] = 2'h0;
    T2[345] = 2'h0;
    T2[346] = 2'h2;
    T2[347] = 2'h1;
    T2[348] = 2'h2;
    T2[349] = 2'h0;
    T2[350] = 2'h1;
    T2[351] = 2'h2;
    T2[352] = 2'h1;
    T2[353] = 2'h2;
    T2[354] = 2'h0;
    T2[355] = 2'h2;
    T2[356] = 2'h2;
    T2[357] = 2'h1;
    T2[358] = 2'h2;
    T2[359] = 2'h0;
    T2[360] = 2'h0;
    T2[361] = 2'h0;
    T2[362] = 2'h2;
    T2[363] = 2'h2;
    T2[364] = 2'h0;
    T2[365] = 2'h1;
    T2[366] = 2'h0;
    T2[367] = 2'h2;
    T2[368] = 2'h2;
    T2[369] = 2'h0;
    T2[370] = 2'h2;
    T2[371] = 2'h0;
    T2[372] = 2'h2;
    T2[373] = 2'h2;
    T2[374] = 2'h0;
    T2[375] = 2'h0;
    T2[376] = 2'h1;
    T2[377] = 2'h2;
    T2[378] = 2'h2;
    T2[379] = 2'h0;
    T2[380] = 2'h1;
    T2[381] = 2'h1;
    T2[382] = 2'h2;
    T2[383] = 2'h2;
    T2[384] = 2'h0;
    T2[385] = 2'h2;
    T2[386] = 2'h1;
    T2[387] = 2'h2;
    T2[388] = 2'h2;
    T2[389] = 2'h0;
    T2[390] = 2'h0;
    T2[391] = 2'h2;
    T2[392] = 2'h2;
    T2[393] = 2'h2;
    T2[394] = 2'h0;
    T2[395] = 2'h1;
    T2[396] = 2'h2;
    T2[397] = 2'h2;
    T2[398] = 2'h2;
    T2[399] = 2'h0;
    T2[400] = 2'h2;
    T2[401] = 2'h2;
    T2[402] = 2'h2;
    T2[403] = 2'h2;
    T2[404] = 2'h0;
    T2[405] = 2'h0;
    T2[406] = 2'h0;
    T2[407] = 2'h0;
    T2[408] = 2'h0;
    T2[409] = 2'h1;
    T2[410] = 2'h1;
    T2[411] = 2'h0;
    T2[412] = 2'h0;
    T2[413] = 2'h0;
    T2[414] = 2'h1;
    T2[415] = 2'h2;
    T2[416] = 2'h0;
    T2[417] = 2'h0;
    T2[418] = 2'h0;
    T2[419] = 2'h1;
    T2[420] = 2'h0;
    T2[421] = 2'h1;
    T2[422] = 2'h0;
    T2[423] = 2'h0;
    T2[424] = 2'h1;
    T2[425] = 2'h1;
    T2[426] = 2'h1;
    T2[427] = 2'h0;
    T2[428] = 2'h0;
    T2[429] = 2'h1;
    T2[430] = 2'h2;
    T2[431] = 2'h1;
    T2[432] = 2'h0;
    T2[433] = 2'h0;
    T2[434] = 2'h1;
    T2[435] = 2'h0;
    T2[436] = 2'h2;
    T2[437] = 2'h0;
    T2[438] = 2'h0;
    T2[439] = 2'h1;
    T2[440] = 2'h1;
    T2[441] = 2'h2;
    T2[442] = 2'h0;
    T2[443] = 2'h0;
    T2[444] = 2'h1;
    T2[445] = 2'h2;
    T2[446] = 2'h2;
    T2[447] = 2'h0;
    T2[448] = 2'h0;
    T2[449] = 2'h1;
    T2[450] = 2'h0;
    T2[451] = 2'h0;
    T2[452] = 2'h1;
    T2[453] = 2'h0;
    T2[454] = 2'h1;
    T2[455] = 2'h1;
    T2[456] = 2'h0;
    T2[457] = 2'h1;
    T2[458] = 2'h0;
    T2[459] = 2'h1;
    T2[460] = 2'h2;
    T2[461] = 2'h0;
    T2[462] = 2'h1;
    T2[463] = 2'h0;
    T2[464] = 2'h1;
    T2[465] = 2'h0;
    T2[466] = 2'h1;
    T2[467] = 2'h1;
    T2[468] = 2'h0;
    T2[469] = 2'h1;
    T2[470] = 2'h1;
    T2[471] = 2'h1;
    T2[472] = 2'h1;
    T2[473] = 2'h0;
    T2[474] = 2'h1;
    T2[475] = 2'h2;
    T2[476] = 2'h1;
    T2[477] = 2'h1;
    T2[478] = 2'h0;
    T2[479] = 2'h1;
    T2[480] = 2'h0;
    T2[481] = 2'h2;
    T2[482] = 2'h1;
    T2[483] = 2'h0;
    T2[484] = 2'h1;
    T2[485] = 2'h1;
    T2[486] = 2'h2;
    T2[487] = 2'h1;
    T2[488] = 2'h0;
    T2[489] = 2'h1;
    T2[490] = 2'h2;
    T2[491] = 2'h2;
    T2[492] = 2'h1;
    T2[493] = 2'h0;
    T2[494] = 2'h1;
    T2[495] = 2'h0;
    T2[496] = 2'h0;
    T2[497] = 2'h2;
    T2[498] = 2'h0;
    T2[499] = 2'h1;
    T2[500] = 2'h1;
    T2[501] = 2'h0;
    T2[502] = 2'h2;
    T2[503] = 2'h0;
    T2[504] = 2'h1;
    T2[505] = 2'h2;
    T2[506] = 2'h0;
    T2[507] = 2'h2;
    T2[508] = 2'h0;
    T2[509] = 2'h1;
    T2[510] = 2'h0;
    T2[511] = 2'h1;
    T2[512] = 2'h2;
    T2[513] = 2'h0;
    T2[514] = 2'h1;
    T2[515] = 2'h1;
    T2[516] = 2'h1;
    T2[517] = 2'h2;
    T2[518] = 2'h0;
    T2[519] = 2'h1;
    T2[520] = 2'h2;
    T2[521] = 2'h1;
    T2[522] = 2'h2;
    T2[523] = 2'h0;
    T2[524] = 2'h1;
    T2[525] = 2'h0;
    T2[526] = 2'h2;
    T2[527] = 2'h2;
    T2[528] = 2'h0;
    T2[529] = 2'h1;
    T2[530] = 2'h1;
    T2[531] = 2'h2;
    T2[532] = 2'h2;
    T2[533] = 2'h0;
    T2[534] = 2'h1;
    T2[535] = 2'h2;
    T2[536] = 2'h2;
    T2[537] = 2'h2;
    T2[538] = 2'h0;
    T2[539] = 2'h1;
    T2[540] = 2'h0;
    T2[541] = 2'h0;
    T2[542] = 2'h0;
    T2[543] = 2'h1;
    T2[544] = 2'h1;
    T2[545] = 2'h1;
    T2[546] = 2'h0;
    T2[547] = 2'h0;
    T2[548] = 2'h1;
    T2[549] = 2'h1;
    T2[550] = 2'h2;
    T2[551] = 2'h0;
    T2[552] = 2'h0;
    T2[553] = 2'h1;
    T2[554] = 2'h1;
    T2[555] = 2'h0;
    T2[556] = 2'h1;
    T2[557] = 2'h0;
    T2[558] = 2'h1;
    T2[559] = 2'h1;
    T2[560] = 2'h1;
    T2[561] = 2'h1;
    T2[562] = 2'h0;
    T2[563] = 2'h1;
    T2[564] = 2'h1;
    T2[565] = 2'h2;
    T2[566] = 2'h1;
    T2[567] = 2'h0;
    T2[568] = 2'h1;
    T2[569] = 2'h1;
    T2[570] = 2'h0;
    T2[571] = 2'h2;
    T2[572] = 2'h0;
    T2[573] = 2'h1;
    T2[574] = 2'h1;
    T2[575] = 2'h1;
    T2[576] = 2'h2;
    T2[577] = 2'h0;
    T2[578] = 2'h1;
    T2[579] = 2'h1;
    T2[580] = 2'h2;
    T2[581] = 2'h2;
    T2[582] = 2'h0;
    T2[583] = 2'h1;
    T2[584] = 2'h1;
    T2[585] = 2'h0;
    T2[586] = 2'h0;
    T2[587] = 2'h1;
    T2[588] = 2'h1;
    T2[589] = 2'h1;
    T2[590] = 2'h1;
    T2[591] = 2'h0;
    T2[592] = 2'h1;
    T2[593] = 2'h1;
    T2[594] = 2'h1;
    T2[595] = 2'h2;
    T2[596] = 2'h0;
    T2[597] = 2'h1;
    T2[598] = 2'h1;
    T2[599] = 2'h1;
    T2[600] = 2'h0;
    T2[601] = 2'h1;
    T2[602] = 2'h1;
    T2[603] = 2'h1;
    T2[604] = 2'h1;
    T2[605] = 2'h1;
    T2[606] = 2'h1;
    T2[607] = 2'h1;
    T2[608] = 2'h1;
    T2[609] = 2'h1;
    T2[610] = 2'h2;
    T2[611] = 2'h1;
    T2[612] = 2'h1;
    T2[613] = 2'h1;
    T2[614] = 2'h1;
    T2[615] = 2'h0;
    T2[616] = 2'h2;
    T2[617] = 2'h1;
    T2[618] = 2'h1;
    T2[619] = 2'h1;
    T2[620] = 2'h1;
    T2[621] = 2'h2;
    T2[622] = 2'h1;
    T2[623] = 2'h1;
    T2[624] = 2'h1;
    T2[625] = 2'h2;
    T2[626] = 2'h2;
    T2[627] = 2'h1;
    T2[628] = 2'h1;
    T2[629] = 2'h1;
    T2[630] = 2'h0;
    T2[631] = 2'h0;
    T2[632] = 2'h2;
    T2[633] = 2'h1;
    T2[634] = 2'h1;
    T2[635] = 2'h1;
    T2[636] = 2'h0;
    T2[637] = 2'h2;
    T2[638] = 2'h1;
    T2[639] = 2'h1;
    T2[640] = 2'h2;
    T2[641] = 2'h0;
    T2[642] = 2'h2;
    T2[643] = 2'h1;
    T2[644] = 2'h1;
    T2[645] = 2'h0;
    T2[646] = 2'h1;
    T2[647] = 2'h2;
    T2[648] = 2'h1;
    T2[649] = 2'h1;
    T2[650] = 2'h1;
    T2[651] = 2'h1;
    T2[652] = 2'h2;
    T2[653] = 2'h1;
    T2[654] = 2'h1;
    T2[655] = 2'h2;
    T2[656] = 2'h1;
    T2[657] = 2'h2;
    T2[658] = 2'h1;
    T2[659] = 2'h1;
    T2[660] = 2'h0;
    T2[661] = 2'h2;
    T2[662] = 2'h2;
    T2[663] = 2'h1;
    T2[664] = 2'h1;
    T2[665] = 2'h1;
    T2[666] = 2'h2;
    T2[667] = 2'h2;
    T2[668] = 2'h1;
    T2[669] = 2'h1;
    T2[670] = 2'h2;
    T2[671] = 2'h2;
    T2[672] = 2'h2;
    T2[673] = 2'h1;
    T2[674] = 2'h1;
    T2[675] = 2'h0;
    T2[676] = 2'h0;
    T2[677] = 2'h0;
    T2[678] = 2'h2;
    T2[679] = 2'h1;
    T2[680] = 2'h1;
    T2[681] = 2'h0;
    T2[682] = 2'h0;
    T2[683] = 2'h2;
    T2[684] = 2'h1;
    T2[685] = 2'h2;
    T2[686] = 2'h0;
    T2[687] = 2'h0;
    T2[688] = 2'h2;
    T2[689] = 2'h1;
    T2[690] = 2'h0;
    T2[691] = 2'h1;
    T2[692] = 2'h0;
    T2[693] = 2'h2;
    T2[694] = 2'h1;
    T2[695] = 2'h1;
    T2[696] = 2'h1;
    T2[697] = 2'h0;
    T2[698] = 2'h2;
    T2[699] = 2'h1;
    T2[700] = 2'h2;
    T2[701] = 2'h1;
    T2[702] = 2'h0;
    T2[703] = 2'h2;
    T2[704] = 2'h1;
    T2[705] = 2'h0;
    T2[706] = 2'h2;
    T2[707] = 2'h0;
    T2[708] = 2'h2;
    T2[709] = 2'h1;
    T2[710] = 2'h1;
    T2[711] = 2'h2;
    T2[712] = 2'h0;
    T2[713] = 2'h2;
    T2[714] = 2'h1;
    T2[715] = 2'h2;
    T2[716] = 2'h2;
    T2[717] = 2'h0;
    T2[718] = 2'h2;
    T2[719] = 2'h1;
    T2[720] = 2'h0;
    T2[721] = 2'h0;
    T2[722] = 2'h1;
    T2[723] = 2'h2;
    T2[724] = 2'h1;
    T2[725] = 2'h1;
    T2[726] = 2'h0;
    T2[727] = 2'h1;
    T2[728] = 2'h2;
    T2[729] = 2'h1;
    T2[730] = 2'h2;
    T2[731] = 2'h0;
    T2[732] = 2'h1;
    T2[733] = 2'h2;
    T2[734] = 2'h1;
    T2[735] = 2'h0;
    T2[736] = 2'h1;
    T2[737] = 2'h1;
    T2[738] = 2'h2;
    T2[739] = 2'h1;
    T2[740] = 2'h1;
    T2[741] = 2'h1;
    T2[742] = 2'h1;
    T2[743] = 2'h2;
    T2[744] = 2'h1;
    T2[745] = 2'h2;
    T2[746] = 2'h1;
    T2[747] = 2'h1;
    T2[748] = 2'h2;
    T2[749] = 2'h1;
    T2[750] = 2'h0;
    T2[751] = 2'h2;
    T2[752] = 2'h1;
    T2[753] = 2'h2;
    T2[754] = 2'h1;
    T2[755] = 2'h1;
    T2[756] = 2'h2;
    T2[757] = 2'h1;
    T2[758] = 2'h2;
    T2[759] = 2'h1;
    T2[760] = 2'h2;
    T2[761] = 2'h2;
    T2[762] = 2'h1;
    T2[763] = 2'h2;
    T2[764] = 2'h1;
    T2[765] = 2'h0;
    T2[766] = 2'h0;
    T2[767] = 2'h2;
    T2[768] = 2'h2;
    T2[769] = 2'h1;
    T2[770] = 2'h1;
    T2[771] = 2'h0;
    T2[772] = 2'h2;
    T2[773] = 2'h2;
    T2[774] = 2'h1;
    T2[775] = 2'h2;
    T2[776] = 2'h0;
    T2[777] = 2'h2;
    T2[778] = 2'h2;
    T2[779] = 2'h1;
    T2[780] = 2'h0;
    T2[781] = 2'h1;
    T2[782] = 2'h2;
    T2[783] = 2'h2;
    T2[784] = 2'h1;
    T2[785] = 2'h1;
    T2[786] = 2'h1;
    T2[787] = 2'h2;
    T2[788] = 2'h2;
    T2[789] = 2'h1;
    T2[790] = 2'h2;
    T2[791] = 2'h1;
    T2[792] = 2'h2;
    T2[793] = 2'h2;
    T2[794] = 2'h1;
    T2[795] = 2'h0;
    T2[796] = 2'h2;
    T2[797] = 2'h2;
    T2[798] = 2'h2;
    T2[799] = 2'h1;
    T2[800] = 2'h1;
    T2[801] = 2'h2;
    T2[802] = 2'h2;
    T2[803] = 2'h2;
    T2[804] = 2'h1;
    T2[805] = 2'h2;
    T2[806] = 2'h2;
    T2[807] = 2'h2;
    T2[808] = 2'h2;
    T2[809] = 2'h1;
    T2[810] = 2'h0;
    T2[811] = 2'h0;
    T2[812] = 2'h0;
    T2[813] = 2'h0;
    T2[814] = 2'h2;
    T2[815] = 2'h1;
    T2[816] = 2'h0;
    T2[817] = 2'h0;
    T2[818] = 2'h0;
    T2[819] = 2'h2;
    T2[820] = 2'h2;
    T2[821] = 2'h0;
    T2[822] = 2'h0;
    T2[823] = 2'h0;
    T2[824] = 2'h2;
    T2[825] = 2'h0;
    T2[826] = 2'h1;
    T2[827] = 2'h0;
    T2[828] = 2'h0;
    T2[829] = 2'h2;
    T2[830] = 2'h1;
    T2[831] = 2'h1;
    T2[832] = 2'h0;
    T2[833] = 2'h0;
    T2[834] = 2'h2;
    T2[835] = 2'h2;
    T2[836] = 2'h1;
    T2[837] = 2'h0;
    T2[838] = 2'h0;
    T2[839] = 2'h2;
    T2[840] = 2'h0;
    T2[841] = 2'h2;
    T2[842] = 2'h0;
    T2[843] = 2'h0;
    T2[844] = 2'h2;
    T2[845] = 2'h1;
    T2[846] = 2'h2;
    T2[847] = 2'h0;
    T2[848] = 2'h0;
    T2[849] = 2'h2;
    T2[850] = 2'h2;
    T2[851] = 2'h2;
    T2[852] = 2'h0;
    T2[853] = 2'h0;
    T2[854] = 2'h2;
    T2[855] = 2'h0;
    T2[856] = 2'h0;
    T2[857] = 2'h1;
    T2[858] = 2'h0;
    T2[859] = 2'h2;
    T2[860] = 2'h1;
    T2[861] = 2'h0;
    T2[862] = 2'h1;
    T2[863] = 2'h0;
    T2[864] = 2'h2;
    T2[865] = 2'h2;
    T2[866] = 2'h0;
    T2[867] = 2'h1;
    T2[868] = 2'h0;
    T2[869] = 2'h2;
    T2[870] = 2'h0;
    T2[871] = 2'h1;
    T2[872] = 2'h1;
    T2[873] = 2'h0;
    T2[874] = 2'h2;
    T2[875] = 2'h1;
    T2[876] = 2'h1;
    T2[877] = 2'h1;
    T2[878] = 2'h0;
    T2[879] = 2'h2;
    T2[880] = 2'h2;
    T2[881] = 2'h1;
    T2[882] = 2'h1;
    T2[883] = 2'h0;
    T2[884] = 2'h2;
    T2[885] = 2'h0;
    T2[886] = 2'h2;
    T2[887] = 2'h1;
    T2[888] = 2'h0;
    T2[889] = 2'h2;
    T2[890] = 2'h1;
    T2[891] = 2'h2;
    T2[892] = 2'h1;
    T2[893] = 2'h0;
    T2[894] = 2'h2;
    T2[895] = 2'h2;
    T2[896] = 2'h2;
    T2[897] = 2'h1;
    T2[898] = 2'h0;
    T2[899] = 2'h2;
    T2[900] = 2'h0;
    T2[901] = 2'h0;
    T2[902] = 2'h2;
    T2[903] = 2'h0;
    T2[904] = 2'h2;
    T2[905] = 2'h1;
    T2[906] = 2'h0;
    T2[907] = 2'h2;
    T2[908] = 2'h0;
    T2[909] = 2'h2;
    T2[910] = 2'h2;
    T2[911] = 2'h0;
    T2[912] = 2'h2;
    T2[913] = 2'h0;
    T2[914] = 2'h2;
    T2[915] = 2'h0;
    T2[916] = 2'h1;
    T2[917] = 2'h2;
    T2[918] = 2'h0;
    T2[919] = 2'h2;
    T2[920] = 2'h1;
    T2[921] = 2'h1;
    T2[922] = 2'h2;
    T2[923] = 2'h0;
    T2[924] = 2'h2;
    T2[925] = 2'h2;
    T2[926] = 2'h1;
    T2[927] = 2'h2;
    T2[928] = 2'h0;
    T2[929] = 2'h2;
    T2[930] = 2'h0;
    T2[931] = 2'h2;
    T2[932] = 2'h2;
    T2[933] = 2'h0;
    T2[934] = 2'h2;
    T2[935] = 2'h1;
    T2[936] = 2'h2;
    T2[937] = 2'h2;
    T2[938] = 2'h0;
    T2[939] = 2'h2;
    T2[940] = 2'h2;
    T2[941] = 2'h2;
    T2[942] = 2'h2;
    T2[943] = 2'h0;
    T2[944] = 2'h2;
    T2[945] = 2'h0;
    T2[946] = 2'h0;
    T2[947] = 2'h0;
    T2[948] = 2'h1;
    T2[949] = 2'h2;
    T2[950] = 2'h1;
    T2[951] = 2'h0;
    T2[952] = 2'h0;
    T2[953] = 2'h1;
    T2[954] = 2'h2;
    T2[955] = 2'h2;
    T2[956] = 2'h0;
    T2[957] = 2'h0;
    T2[958] = 2'h1;
    T2[959] = 2'h2;
    T2[960] = 2'h0;
    T2[961] = 2'h1;
    T2[962] = 2'h0;
    T2[963] = 2'h1;
    T2[964] = 2'h2;
    T2[965] = 2'h1;
    T2[966] = 2'h1;
    T2[967] = 2'h0;
    T2[968] = 2'h1;
    T2[969] = 2'h2;
    T2[970] = 2'h2;
    T2[971] = 2'h1;
    T2[972] = 2'h0;
    T2[973] = 2'h1;
    T2[974] = 2'h2;
    T2[975] = 2'h0;
    T2[976] = 2'h2;
    T2[977] = 2'h0;
    T2[978] = 2'h1;
    T2[979] = 2'h2;
    T2[980] = 2'h1;
    T2[981] = 2'h2;
    T2[982] = 2'h0;
    T2[983] = 2'h1;
    T2[984] = 2'h2;
    T2[985] = 2'h2;
    T2[986] = 2'h2;
    T2[987] = 2'h0;
    T2[988] = 2'h1;
    T2[989] = 2'h2;
    T2[990] = 2'h0;
    T2[991] = 2'h0;
    T2[992] = 2'h1;
    T2[993] = 2'h1;
    T2[994] = 2'h2;
    T2[995] = 2'h1;
    T2[996] = 2'h0;
    T2[997] = 2'h1;
    T2[998] = 2'h1;
    T2[999] = 2'h2;
    T2[1000] = 2'h2;
    T2[1001] = 2'h0;
    T2[1002] = 2'h1;
    T2[1003] = 2'h1;
    T2[1004] = 2'h2;
    T2[1005] = 2'h0;
    T2[1006] = 2'h1;
    T2[1007] = 2'h1;
    T2[1008] = 2'h1;
    T2[1009] = 2'h2;
    T2[1010] = 2'h1;
    T2[1011] = 2'h1;
    T2[1012] = 2'h1;
    T2[1013] = 2'h1;
    T2[1014] = 2'h2;
    T2[1015] = 2'h2;
    T2[1016] = 2'h1;
    T2[1017] = 2'h1;
    T2[1018] = 2'h1;
    T2[1019] = 2'h2;
    T2[1020] = 2'h0;
    T2[1021] = 2'h2;
    T2[1022] = 2'h1;
    T2[1023] = 2'h1;
    T2[1024] = 2'h2;
    T2[1025] = 2'h1;
    T2[1026] = 2'h2;
    T2[1027] = 2'h1;
    T2[1028] = 2'h1;
    T2[1029] = 2'h2;
    T2[1030] = 2'h2;
    T2[1031] = 2'h2;
    T2[1032] = 2'h1;
    T2[1033] = 2'h1;
    T2[1034] = 2'h2;
    T2[1035] = 2'h0;
    T2[1036] = 2'h0;
    T2[1037] = 2'h2;
    T2[1038] = 2'h1;
    T2[1039] = 2'h2;
    T2[1040] = 2'h1;
    T2[1041] = 2'h0;
    T2[1042] = 2'h2;
    T2[1043] = 2'h1;
    T2[1044] = 2'h2;
    T2[1045] = 2'h2;
    T2[1046] = 2'h0;
    T2[1047] = 2'h2;
    T2[1048] = 2'h1;
    T2[1049] = 2'h2;
    T2[1050] = 2'h0;
    T2[1051] = 2'h1;
    T2[1052] = 2'h2;
    T2[1053] = 2'h1;
    T2[1054] = 2'h2;
    T2[1055] = 2'h1;
    T2[1056] = 2'h1;
    T2[1057] = 2'h2;
    T2[1058] = 2'h1;
    T2[1059] = 2'h2;
    T2[1060] = 2'h2;
    T2[1061] = 2'h1;
    T2[1062] = 2'h2;
    T2[1063] = 2'h1;
    T2[1064] = 2'h2;
    T2[1065] = 2'h0;
    T2[1066] = 2'h2;
    T2[1067] = 2'h2;
    T2[1068] = 2'h1;
    T2[1069] = 2'h2;
    T2[1070] = 2'h1;
    T2[1071] = 2'h2;
    T2[1072] = 2'h2;
    T2[1073] = 2'h1;
    T2[1074] = 2'h2;
    T2[1075] = 2'h2;
    T2[1076] = 2'h2;
    T2[1077] = 2'h2;
    T2[1078] = 2'h1;
    T2[1079] = 2'h2;
    T2[1080] = 2'h0;
    T2[1081] = 2'h0;
    T2[1082] = 2'h0;
    T2[1083] = 2'h2;
    T2[1084] = 2'h2;
    T2[1085] = 2'h1;
    T2[1086] = 2'h0;
    T2[1087] = 2'h0;
    T2[1088] = 2'h2;
    T2[1089] = 2'h2;
    T2[1090] = 2'h2;
    T2[1091] = 2'h0;
    T2[1092] = 2'h0;
    T2[1093] = 2'h2;
    T2[1094] = 2'h2;
    T2[1095] = 2'h0;
    T2[1096] = 2'h1;
    T2[1097] = 2'h0;
    T2[1098] = 2'h2;
    T2[1099] = 2'h2;
    T2[1100] = 2'h1;
    T2[1101] = 2'h1;
    T2[1102] = 2'h0;
    T2[1103] = 2'h2;
    T2[1104] = 2'h2;
    T2[1105] = 2'h2;
    T2[1106] = 2'h1;
    T2[1107] = 2'h0;
    T2[1108] = 2'h2;
    T2[1109] = 2'h2;
    T2[1110] = 2'h0;
    T2[1111] = 2'h2;
    T2[1112] = 2'h0;
    T2[1113] = 2'h2;
    T2[1114] = 2'h2;
    T2[1115] = 2'h1;
    T2[1116] = 2'h2;
    T2[1117] = 2'h0;
    T2[1118] = 2'h2;
    T2[1119] = 2'h2;
    T2[1120] = 2'h2;
    T2[1121] = 2'h2;
    T2[1122] = 2'h0;
    T2[1123] = 2'h2;
    T2[1124] = 2'h2;
    T2[1125] = 2'h0;
    T2[1126] = 2'h0;
    T2[1127] = 2'h1;
    T2[1128] = 2'h2;
    T2[1129] = 2'h2;
    T2[1130] = 2'h1;
    T2[1131] = 2'h0;
    T2[1132] = 2'h1;
    T2[1133] = 2'h2;
    T2[1134] = 2'h2;
    T2[1135] = 2'h2;
    T2[1136] = 2'h0;
    T2[1137] = 2'h1;
    T2[1138] = 2'h2;
    T2[1139] = 2'h2;
    T2[1140] = 2'h0;
    T2[1141] = 2'h1;
    T2[1142] = 2'h1;
    T2[1143] = 2'h2;
    T2[1144] = 2'h2;
    T2[1145] = 2'h1;
    T2[1146] = 2'h1;
    T2[1147] = 2'h1;
    T2[1148] = 2'h2;
    T2[1149] = 2'h2;
    T2[1150] = 2'h2;
    T2[1151] = 2'h1;
    T2[1152] = 2'h1;
    T2[1153] = 2'h2;
    T2[1154] = 2'h2;
    T2[1155] = 2'h0;
    T2[1156] = 2'h2;
    T2[1157] = 2'h1;
    T2[1158] = 2'h2;
    T2[1159] = 2'h2;
    T2[1160] = 2'h1;
    T2[1161] = 2'h2;
    T2[1162] = 2'h1;
    T2[1163] = 2'h2;
    T2[1164] = 2'h2;
    T2[1165] = 2'h2;
    T2[1166] = 2'h2;
    T2[1167] = 2'h1;
    T2[1168] = 2'h2;
    T2[1169] = 2'h2;
    T2[1170] = 2'h0;
    T2[1171] = 2'h0;
    T2[1172] = 2'h2;
    T2[1173] = 2'h2;
    T2[1174] = 2'h2;
    T2[1175] = 2'h1;
    T2[1176] = 2'h0;
    T2[1177] = 2'h2;
    T2[1178] = 2'h2;
    T2[1179] = 2'h2;
    T2[1180] = 2'h2;
    T2[1181] = 2'h0;
    T2[1182] = 2'h2;
    T2[1183] = 2'h2;
    T2[1184] = 2'h2;
    T2[1185] = 2'h0;
    T2[1186] = 2'h1;
    T2[1187] = 2'h2;
    T2[1188] = 2'h2;
    T2[1189] = 2'h2;
    T2[1190] = 2'h1;
    T2[1191] = 2'h1;
    T2[1192] = 2'h2;
    T2[1193] = 2'h2;
    T2[1194] = 2'h2;
    T2[1195] = 2'h2;
    T2[1196] = 2'h1;
    T2[1197] = 2'h2;
    T2[1198] = 2'h2;
    T2[1199] = 2'h2;
    T2[1200] = 2'h0;
    T2[1201] = 2'h2;
    T2[1202] = 2'h2;
    T2[1203] = 2'h2;
    T2[1204] = 2'h2;
    T2[1205] = 2'h1;
    T2[1206] = 2'h2;
    T2[1207] = 2'h2;
    T2[1208] = 2'h2;
    T2[1209] = 2'h2;
    T2[1210] = 2'h2;
    T2[1211] = 2'h2;
    T2[1212] = 2'h2;
    T2[1213] = 2'h2;
    T2[1214] = 2'h2;
  end
  assign T3 = T4[4'ha:1'h0];
  assign T4 = index + T5;
  assign T5 = {11'h0, io_inb};
  assign index = io_ina * 3'h5;
endmodule

