module radix2345(
    input [3:0] io_radix,
    input [15:0] io_x0_real,
    input [15:0] io_x0_imag,
    input [15:0] io_x1_real,
    input [15:0] io_x1_imag,
    input [15:0] io_x2_real,
    input [15:0] io_x2_imag,
    input [15:0] io_x3_real,
    input [15:0] io_x3_imag,
    input [15:0] io_x4_real,
    input [15:0] io_x4_imag,
    input [15:0] io_twiddle1_real,
    input [15:0] io_twiddle1_imag,
    input [15:0] io_twiddle2_real,
    input [15:0] io_twiddle2_imag,
    input [15:0] io_twiddle3_real,
    input [15:0] io_twiddle3_imag,
    input [15:0] io_twiddle4_real,
    input [15:0] io_twiddle4_imag,
    output[15:0] io_y0_real,
    output[15:0] io_y0_imag,
    output[15:0] io_y1_real,
    output[15:0] io_y1_imag,
    output[15:0] io_y2_real,
    output[15:0] io_y2_imag,
    output[15:0] io_y3_real,
    output[15:0] io_y3_imag,
    output[15:0] io_y4_real,
    output[15:0] io_y4_imag
);

  wire[15:0] T0;
  wire[52:0] T1;
  wire[52:0] T2;
  wire[52:0] T3;
  wire[36:0] T4;
  wire T5;
  wire[52:0] yx4_imag;
  wire[52:0] T6;
  wire[36:0] T7;
  wire[36:0] yz4_real;
  wire[36:0] T8;
  wire[31:0] T9;
  wire[31:0] T10;
  wire[15:0] d4_imag;
  wire[15:0] d42_imag;
  wire[15:0] T11;
  wire[36:0] T12;
  wire[36:0] T13;
  wire[36:0] c6_imag;
  wire[36:0] T14;
  wire[15:0] b6_imag;
  wire[15:0] b4_imag;
  wire[15:0] a42_imag;
  wire[15:0] T15;
  wire[15:0] T16;
  wire[15:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[15:0] b3_imag;
  wire[15:0] a32_imag;
  wire[15:0] T24;
  wire[15:0] T25;
  wire T26;
  wire T27;
  wire[15:0] a31_imag;
  wire[15:0] T28;
  wire[15:0] T29;
  wire T30;
  wire T31;
  wire[15:0] c4_imag;
  wire[15:0] T32;
  wire[36:0] T33;
  wire[36:0] T34;
  wire[36:0] T35;
  wire[35:0] T36;
  wire[35:0] T37;
  wire T38;
  wire[36:0] T39;
  wire[36:0] T40;
  wire[36:0] T41;
  wire T42;
  wire[31:0] T43;
  wire[15:0] T44;
  wire[15:0] d4_real;
  wire[15:0] d42_real;
  wire[15:0] T45;
  wire[36:0] T46;
  wire[36:0] T47;
  wire[36:0] c6_real;
  wire[36:0] T48;
  wire[15:0] b6_real;
  wire[15:0] b4_real;
  wire[15:0] a42_real;
  wire[15:0] T49;
  wire[15:0] T50;
  wire[15:0] T51;
  wire[15:0] b3_real;
  wire[15:0] a32_real;
  wire[15:0] T52;
  wire[15:0] T53;
  wire[15:0] a31_real;
  wire[15:0] T54;
  wire[15:0] T55;
  wire[15:0] c4_real;
  wire[15:0] T56;
  wire[36:0] T57;
  wire[36:0] T58;
  wire[36:0] T59;
  wire[35:0] T60;
  wire[35:0] T61;
  wire T62;
  wire[36:0] T63;
  wire[36:0] T64;
  wire[36:0] T65;
  wire T66;
  wire[4:0] T67;
  wire T68;
  wire[36:0] d1_real;
  wire[36:0] T69;
  wire[15:0] d12_real;
  wire[15:0] T70;
  wire[36:0] T71;
  wire[36:0] T72;
  wire[36:0] c5_real;
  wire[36:0] T73;
  wire[15:0] b5_real;
  wire[15:0] b52_real;
  wire[15:0] T74;
  wire[15:0] T75;
  wire[15:0] b2_real;
  wire[15:0] a22_real;
  wire[15:0] T76;
  wire[15:0] T77;
  wire[15:0] b1_real;
  wire[15:0] a12_real;
  wire[15:0] T78;
  wire[15:0] T79;
  wire[15:0] T80;
  wire[15:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[15:0] b51_real;
  wire[15:0] T92;
  wire[15:0] T93;
  wire[20:0] T94;
  wire T95;
  wire[36:0] c1_real;
  wire[36:0] T96;
  wire[36:0] T97;
  wire[36:0] T98;
  wire[20:0] T99;
  wire T100;
  wire[36:0] yz4_imag;
  wire[36:0] T101;
  wire[31:0] T102;
  wire[31:0] T103;
  wire[4:0] T104;
  wire T105;
  wire[36:0] d1_imag;
  wire[36:0] T106;
  wire[15:0] d12_imag;
  wire[15:0] T107;
  wire[36:0] T108;
  wire[36:0] T109;
  wire[36:0] c5_imag;
  wire[36:0] T110;
  wire[15:0] b5_imag;
  wire[15:0] b52_imag;
  wire[15:0] T111;
  wire[15:0] T112;
  wire[15:0] b2_imag;
  wire[15:0] a22_imag;
  wire[15:0] T113;
  wire[15:0] T114;
  wire[15:0] b1_imag;
  wire[15:0] a12_imag;
  wire[15:0] T115;
  wire[15:0] T116;
  wire[15:0] T117;
  wire[15:0] T118;
  wire[15:0] b51_imag;
  wire[15:0] T119;
  wire[15:0] T120;
  wire[20:0] T121;
  wire T122;
  wire[36:0] c1_imag;
  wire[36:0] T123;
  wire[36:0] T124;
  wire[36:0] T125;
  wire[20:0] T126;
  wire T127;
  wire[52:0] T128;
  wire[15:0] T129;
  wire T130;
  wire[52:0] T131;
  wire[36:0] T132;
  wire T133;
  wire T134;
  wire[15:0] T135;
  wire[52:0] T136;
  wire[52:0] T137;
  wire[52:0] T138;
  wire[36:0] T139;
  wire T140;
  wire[52:0] yx4_real;
  wire[52:0] T141;
  wire[36:0] T142;
  wire[52:0] T143;
  wire[36:0] T144;
  wire T145;
  wire[15:0] T146;
  wire[31:0] T147;
  wire[31:0] T148;
  wire[31:0] T149;
  wire[15:0] T150;
  wire T151;
  wire[31:0] yx3_imag;
  wire[31:0] T152;
  wire[15:0] T153;
  wire[15:0] yy3_real;
  wire[15:0] T154;
  wire[31:0] T155;
  wire[31:0] T156;
  wire[31:0] yz3_real;
  wire[31:0] T157;
  wire[31:0] T158;
  wire[15:0] yz22_imag;
  wire[15:0] T159;
  wire[37:0] T160;
  wire[37:0] T161;
  wire[37:0] d3_imag;
  wire[37:0] T162;
  wire T163;
  wire[37:0] c3_imag;
  wire[37:0] T164;
  wire[37:0] T165;
  wire[21:0] T166;
  wire T167;
  wire[31:0] T168;
  wire[15:0] T169;
  wire[15:0] yz22_real;
  wire[15:0] T170;
  wire[37:0] T171;
  wire[37:0] T172;
  wire[37:0] d3_real;
  wire[37:0] T173;
  wire T174;
  wire[37:0] c3_real;
  wire[37:0] T175;
  wire[37:0] T176;
  wire[21:0] T177;
  wire T178;
  wire[31:0] T179;
  wire[15:0] yz21_real;
  wire[15:0] T180;
  wire[36:0] T181;
  wire[36:0] T182;
  wire[36:0] d2_real;
  wire[36:0] T183;
  wire[15:0] c2_real;
  wire[15:0] c22_real;
  wire[15:0] T184;
  wire[36:0] T185;
  wire[36:0] T186;
  wire[36:0] T187;
  wire[36:0] T188;
  wire[36:0] T189;
  wire[20:0] T190;
  wire T191;
  wire T192;
  wire T193;
  wire[20:0] T194;
  wire T195;
  wire[36:0] T196;
  wire[20:0] T197;
  wire T198;
  wire[15:0] T199;
  wire T200;
  wire[31:0] yz2_real;
  wire[31:0] T201;
  wire[31:0] T202;
  wire[31:0] T203;
  wire[15:0] T204;
  wire[31:0] T205;
  wire[15:0] T206;
  wire T207;
  wire[15:0] yy3_imag;
  wire[15:0] T208;
  wire[31:0] T209;
  wire[31:0] T210;
  wire[31:0] yz3_imag;
  wire[31:0] T211;
  wire[31:0] T212;
  wire[31:0] T213;
  wire[15:0] yz21_imag;
  wire[15:0] T214;
  wire[36:0] T215;
  wire[36:0] T216;
  wire[36:0] d2_imag;
  wire[36:0] T217;
  wire[15:0] c2_imag;
  wire[15:0] c22_imag;
  wire[15:0] T218;
  wire[36:0] T219;
  wire[36:0] T220;
  wire[36:0] T221;
  wire[36:0] T222;
  wire[36:0] T223;
  wire[20:0] T224;
  wire T225;
  wire[20:0] T226;
  wire T227;
  wire[36:0] T228;
  wire[20:0] T229;
  wire T230;
  wire[15:0] T231;
  wire T232;
  wire[31:0] yz2_imag;
  wire[31:0] T233;
  wire[31:0] T234;
  wire[31:0] T235;
  wire[15:0] T236;
  wire T237;
  wire[31:0] T238;
  wire[15:0] T239;
  wire T240;
  wire[31:0] T241;
  wire[15:0] T242;
  wire T243;
  wire T244;
  wire[15:0] T245;
  wire[31:0] T246;
  wire[31:0] T247;
  wire[31:0] T248;
  wire[15:0] T249;
  wire T250;
  wire[31:0] yx3_real;
  wire[31:0] T251;
  wire[15:0] T252;
  wire[31:0] T253;
  wire[15:0] T254;
  wire T255;
  wire[15:0] T256;
  wire[31:0] T257;
  wire[31:0] T258;
  wire[31:0] T259;
  wire[15:0] T260;
  wire T261;
  wire[31:0] yx2_imag;
  wire[31:0] T262;
  wire[15:0] T263;
  wire[15:0] yy2_real;
  wire[15:0] T264;
  wire[36:0] T265;
  wire[36:0] T266;
  wire[36:0] T267;
  wire[36:0] T268;
  wire[4:0] T269;
  wire T270;
  wire[36:0] T271;
  wire[20:0] T272;
  wire T273;
  wire[36:0] T274;
  wire[4:0] T275;
  wire T276;
  wire[15:0] yy2_imag;
  wire[15:0] T277;
  wire[36:0] T278;
  wire[36:0] T279;
  wire[36:0] T280;
  wire[36:0] T281;
  wire[4:0] T282;
  wire T283;
  wire[36:0] T284;
  wire[20:0] T285;
  wire T286;
  wire[36:0] T287;
  wire[4:0] T288;
  wire T289;
  wire[31:0] T290;
  wire[15:0] T291;
  wire T292;
  wire[31:0] T293;
  wire[15:0] T294;
  wire T295;
  wire T296;
  wire[15:0] T297;
  wire[31:0] T298;
  wire[31:0] T299;
  wire[31:0] T300;
  wire[15:0] T301;
  wire T302;
  wire[31:0] yx2_real;
  wire[31:0] T303;
  wire[15:0] T304;
  wire[31:0] T305;
  wire[15:0] T306;
  wire T307;
  wire[15:0] T308;
  wire[31:0] T309;
  wire[31:0] T310;
  wire[15:0] T311;
  wire[15:0] yy1_real;
  wire[15:0] T312;
  wire[36:0] T313;
  wire[36:0] T314;
  wire[36:0] T315;
  wire[36:0] T316;
  wire[36:0] yz1_real;
  wire[36:0] T317;
  wire[31:0] T318;
  wire[31:0] T319;
  wire[31:0] T320;
  wire[15:0] T321;
  wire[4:0] T322;
  wire T323;
  wire[36:0] T324;
  wire[20:0] T325;
  wire T326;
  wire[36:0] T327;
  wire[4:0] T328;
  wire T329;
  wire[15:0] yy1_imag;
  wire[15:0] T330;
  wire[36:0] T331;
  wire[36:0] T332;
  wire[36:0] T333;
  wire[36:0] T334;
  wire[36:0] yz1_imag;
  wire[36:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[4:0] T338;
  wire T339;
  wire[36:0] T340;
  wire[20:0] T341;
  wire T342;
  wire[36:0] T343;
  wire[4:0] T344;
  wire T345;
  wire[31:0] T346;
  wire[15:0] T347;
  wire[15:0] T348;
  wire[31:0] T349;
  wire[31:0] T350;
  wire[15:0] T351;
  wire[15:0] T352;
  wire[15:0] T353;
  wire[15:0] T354;
  wire[15:0] T355;
  wire[15:0] yz0_imag;
  wire[15:0] d02_imag;
  wire[15:0] T356;
  wire[15:0] T357;
  wire[15:0] c7_imag;
  wire[15:0] T358;
  wire[15:0] T359;
  wire[15:0] T360;
  wire[15:0] T361;
  wire[15:0] yz0_real;
  wire[15:0] d02_real;
  wire[15:0] T362;
  wire[15:0] T363;
  wire[15:0] c7_real;


  assign io_y4_imag = T0;
  assign T0 = T1[4'hf:1'h0];
  assign T1 = T134 ? T131 : T2;
  assign T2 = T130 ? yx4_imag : T3;
  assign T3 = {T4, io_x4_imag};
  assign T4 = T5 ? 37'h1fffffffff : 37'h0;
  assign T5 = io_x4_imag[4'hf:4'hf];
  assign yx4_imag = T128 + T6;
  assign T6 = $signed(T7) * $signed(io_twiddle4_real);
  assign T7 = yz4_imag - yz4_real;
  assign yz4_real = d1_real - T8;
  assign T8 = {T67, T9};
  assign T9 = T43 - T10;
  assign T10 = $signed(16'h1) * $signed(d4_imag);
  assign d4_imag = c4_imag + d42_imag;
  assign d42_imag = T11;
  assign T11 = T12[4'hf:1'h0];
  assign T12 = T31 ? c6_imag : T13;
  assign T13 = T30 ? 37'h0 : c6_imag;
  assign c6_imag = $signed(T14) / $signed(22'h100000);
  assign T14 = $signed(21'h16986f) * $signed(b6_imag);
  assign b6_imag = b3_imag + b4_imag;
  assign b4_imag = io_x1_imag - a42_imag;
  assign a42_imag = T15;
  assign T15 = T22 ? io_x4_imag : T16;
  assign T16 = T19 ? io_x3_imag : T17;
  assign T17 = T18 ? io_x2_imag : io_x4_imag;
  assign T18 = io_radix == 4'h3;
  assign T19 = T21 & T20;
  assign T20 = io_radix == 4'h4;
  assign T21 = T18 == 1'h0;
  assign T22 = T23 == 1'h0;
  assign T23 = T18 | T20;
  assign b3_imag = a31_imag - a32_imag;
  assign a32_imag = T24;
  assign T24 = T27 ? io_x3_imag : T25;
  assign T25 = T26 ? io_x2_imag : io_x3_imag;
  assign T26 = io_radix == 4'h4;
  assign T27 = T26 == 1'h0;
  assign a31_imag = T28;
  assign T28 = T27 ? io_x2_imag : T29;
  assign T29 = T26 ? io_x0_imag : io_x2_imag;
  assign T30 = io_radix == 4'h3;
  assign T31 = T30 == 1'h0;
  assign c4_imag = T32;
  assign T32 = T33[4'hf:1'h0];
  assign T33 = T31 ? T41 : T34;
  assign T34 = T30 ? T39 : T35;
  assign T35 = {T38, T36};
  assign T36 = $signed(T37) / $signed(22'h100000);
  assign T37 = $signed(20'ha300b) * $signed(b4_imag);
  assign T38 = T36[6'h23:6'h23];
  assign T39 = $signed(T40) / $signed(22'h100000);
  assign T40 = $signed(21'h1224c3) * $signed(b4_imag);
  assign T41 = {T42, T36};
  assign T42 = T36[6'h23:6'h23];
  assign T43 = $signed(16'h0) * $signed(T44);
  assign T44 = d4_real + d4_imag;
  assign d4_real = c4_real + d42_real;
  assign d42_real = T45;
  assign T45 = T46[4'hf:1'h0];
  assign T46 = T31 ? c6_real : T47;
  assign T47 = T30 ? 37'h0 : c6_real;
  assign c6_real = $signed(T48) / $signed(22'h100000);
  assign T48 = $signed(21'h16986f) * $signed(b6_real);
  assign b6_real = b3_real + b4_real;
  assign b4_real = io_x1_real - a42_real;
  assign a42_real = T49;
  assign T49 = T22 ? io_x4_real : T50;
  assign T50 = T19 ? io_x3_real : T51;
  assign T51 = T18 ? io_x2_real : io_x4_real;
  assign b3_real = a31_real - a32_real;
  assign a32_real = T52;
  assign T52 = T27 ? io_x3_real : T53;
  assign T53 = T26 ? io_x2_real : io_x3_real;
  assign a31_real = T54;
  assign T54 = T27 ? io_x2_real : T55;
  assign T55 = T26 ? io_x0_real : io_x2_real;
  assign c4_real = T56;
  assign T56 = T57[4'hf:1'h0];
  assign T57 = T31 ? T65 : T58;
  assign T58 = T30 ? T63 : T59;
  assign T59 = {T62, T60};
  assign T60 = $signed(T61) / $signed(22'h100000);
  assign T61 = $signed(20'ha300b) * $signed(b4_real);
  assign T62 = T60[6'h23:6'h23];
  assign T63 = $signed(T64) / $signed(22'h100000);
  assign T64 = $signed(21'h1224c3) * $signed(b4_real);
  assign T65 = {T66, T60};
  assign T66 = T60[6'h23:6'h23];
  assign T67 = T68 ? 5'h1f : 5'h0;
  assign T68 = T9[5'h1f:5'h1f];
  assign d1_real = c1_real - T69;
  assign T69 = {T94, d12_real};
  assign d12_real = T70;
  assign T70 = T71[4'hf:1'h0];
  assign T71 = T31 ? c5_real : T72;
  assign T72 = T30 ? 37'h0 : c5_real;
  assign c5_real = $signed(T73) / $signed(22'h100000);
  assign T73 = $signed(21'h130e45) * $signed(b5_real);
  assign b5_real = b51_real - b52_real;
  assign b52_real = T74;
  assign T74 = T27 ? b2_real : T75;
  assign T75 = T26 ? b1_real : b2_real;
  assign b2_real = io_x2_real + a22_real;
  assign a22_real = T76;
  assign T76 = T27 ? io_x3_real : T77;
  assign T77 = T26 ? io_x0_real : io_x3_real;
  assign b1_real = io_x1_real + a12_real;
  assign a12_real = T78;
  assign T78 = T90 ? io_x4_real : T79;
  assign T79 = T86 ? io_x3_real : T80;
  assign T80 = T83 ? io_x2_real : T81;
  assign T81 = T82 ? io_x0_real : io_x4_real;
  assign T82 = io_radix == 4'h2;
  assign T83 = T85 & T84;
  assign T84 = io_radix == 4'h3;
  assign T85 = T82 == 1'h0;
  assign T86 = T88 & T87;
  assign T87 = io_radix == 4'h4;
  assign T88 = T89 == 1'h0;
  assign T89 = T82 | T84;
  assign T90 = T91 == 1'h0;
  assign T91 = T89 | T87;
  assign b51_real = T92;
  assign T92 = T27 ? b1_real : T93;
  assign T93 = T26 ? b2_real : b1_real;
  assign T94 = T95 ? 21'h1fffff : 21'h0;
  assign T95 = d12_real[4'hf:4'hf];
  assign c1_real = T98 - T96;
  assign T96 = $signed(T97) / $signed(22'h100000);
  assign T97 = $signed(21'h80000) * $signed(b1_real);
  assign T98 = {T99, io_x0_real};
  assign T99 = T100 ? 21'h1fffff : 21'h0;
  assign T100 = io_x0_real[4'hf:4'hf];
  assign yz4_imag = d1_imag - T101;
  assign T101 = {T104, T102};
  assign T102 = T43 + T103;
  assign T103 = $signed(16'h1) * $signed(d4_real);
  assign T104 = T105 ? 5'h1f : 5'h0;
  assign T105 = T102[5'h1f:5'h1f];
  assign d1_imag = c1_imag - T106;
  assign T106 = {T121, d12_imag};
  assign d12_imag = T107;
  assign T107 = T108[4'hf:1'h0];
  assign T108 = T31 ? c5_imag : T109;
  assign T109 = T30 ? 37'h0 : c5_imag;
  assign c5_imag = $signed(T110) / $signed(22'h100000);
  assign T110 = $signed(21'h130e45) * $signed(b5_imag);
  assign b5_imag = b51_imag - b52_imag;
  assign b52_imag = T111;
  assign T111 = T27 ? b2_imag : T112;
  assign T112 = T26 ? b1_imag : b2_imag;
  assign b2_imag = io_x2_imag + a22_imag;
  assign a22_imag = T113;
  assign T113 = T27 ? io_x3_imag : T114;
  assign T114 = T26 ? io_x0_imag : io_x3_imag;
  assign b1_imag = io_x1_imag + a12_imag;
  assign a12_imag = T115;
  assign T115 = T90 ? io_x4_imag : T116;
  assign T116 = T86 ? io_x3_imag : T117;
  assign T117 = T83 ? io_x2_imag : T118;
  assign T118 = T82 ? io_x0_imag : io_x4_imag;
  assign b51_imag = T119;
  assign T119 = T27 ? b1_imag : T120;
  assign T120 = T26 ? b2_imag : b1_imag;
  assign T121 = T122 ? 21'h1fffff : 21'h0;
  assign T122 = d12_imag[4'hf:4'hf];
  assign c1_imag = T125 - T123;
  assign T123 = $signed(T124) / $signed(22'h100000);
  assign T124 = $signed(21'h80000) * $signed(b1_imag);
  assign T125 = {T126, io_x0_imag};
  assign T126 = T127 ? 21'h1fffff : 21'h0;
  assign T127 = io_x0_imag[4'hf:4'hf];
  assign T128 = $signed(yz4_real) * $signed(T129);
  assign T129 = io_twiddle4_real + io_twiddle4_imag;
  assign T130 = 4'h4 < io_radix;
  assign T131 = {T132, io_x4_imag};
  assign T132 = T133 ? 37'h1fffffffff : 37'h0;
  assign T133 = io_x4_imag[4'hf:4'hf];
  assign T134 = T130 == 1'h0;
  assign io_y4_real = T135;
  assign T135 = T136[4'hf:1'h0];
  assign T136 = T134 ? T143 : T137;
  assign T137 = T130 ? yx4_real : T138;
  assign T138 = {T139, io_x4_real};
  assign T139 = T140 ? 37'h1fffffffff : 37'h0;
  assign T140 = io_x4_real[4'hf:4'hf];
  assign yx4_real = T128 - T141;
  assign T141 = $signed(T142) * $signed(io_twiddle4_imag);
  assign T142 = yz4_real + yz4_imag;
  assign T143 = {T144, io_x4_real};
  assign T144 = T145 ? 37'h1fffffffff : 37'h0;
  assign T145 = io_x4_real[4'hf:4'hf];
  assign io_y3_imag = T146;
  assign T146 = T147[4'hf:1'h0];
  assign T147 = T244 ? T241 : T148;
  assign T148 = T240 ? yx3_imag : T149;
  assign T149 = {T150, io_x3_imag};
  assign T150 = T151 ? 16'hffff : 16'h0;
  assign T151 = io_x3_imag[4'hf:4'hf];
  assign yx3_imag = T238 + T152;
  assign T152 = $signed(T153) * $signed(io_twiddle3_real);
  assign T153 = yy3_imag - yy3_real;
  assign yy3_real = T154;
  assign T154 = T155[4'hf:1'h0];
  assign T155 = T27 ? yz3_real : T156;
  assign T156 = T26 ? yz2_real : yz3_real;
  assign yz3_real = T179 - T157;
  assign T157 = T168 - T158;
  assign T158 = $signed(16'h1) * $signed(yz22_imag);
  assign yz22_imag = T159;
  assign T159 = T160[4'hf:1'h0];
  assign T160 = T27 ? d3_imag : T161;
  assign T161 = T26 ? T165 : d3_imag;
  assign d3_imag = c3_imag + T162;
  assign T162 = {T163, c6_imag};
  assign T163 = c6_imag[6'h24:6'h24];
  assign c3_imag = $signed(T164) / $signed(22'h100000);
  assign T164 = $signed(22'h189f18) * $signed(b3_imag);
  assign T165 = {T166, b4_imag};
  assign T166 = T167 ? 22'h3fffff : 22'h0;
  assign T167 = b4_imag[4'hf:4'hf];
  assign T168 = $signed(16'h0) * $signed(T169);
  assign T169 = yz22_real + yz22_imag;
  assign yz22_real = T170;
  assign T170 = T171[4'hf:1'h0];
  assign T171 = T27 ? d3_real : T172;
  assign T172 = T26 ? T176 : d3_real;
  assign d3_real = c3_real + T173;
  assign T173 = {T174, c6_real};
  assign T174 = c6_real[6'h24:6'h24];
  assign c3_real = $signed(T175) / $signed(22'h100000);
  assign T175 = $signed(22'h189f18) * $signed(b3_real);
  assign T176 = {T177, b4_real};
  assign T177 = T178 ? 22'h3fffff : 22'h0;
  assign T178 = b4_real[4'hf:4'hf];
  assign T179 = {T199, yz21_real};
  assign yz21_real = T180;
  assign T180 = T181[4'hf:1'h0];
  assign T181 = T27 ? d2_real : T182;
  assign T182 = T26 ? T196 : d2_real;
  assign d2_real = T183 + c5_real;
  assign T183 = {T194, c2_real};
  assign c2_real = io_x0_real - c22_real;
  assign c22_real = T184;
  assign T184 = T185[4'hf:1'h0];
  assign T185 = T193 ? T187 : T186;
  assign T186 = T192 ? T189 : T187;
  assign T187 = $signed(T188) / $signed(22'h100000);
  assign T188 = $signed(21'h80000) * $signed(b2_real);
  assign T189 = {T190, io_x1_real};
  assign T190 = T191 ? 21'h1fffff : 21'h0;
  assign T191 = io_x1_real[4'hf:4'hf];
  assign T192 = io_radix == 4'h2;
  assign T193 = T192 == 1'h0;
  assign T194 = T195 ? 21'h1fffff : 21'h0;
  assign T195 = c2_real[4'hf:4'hf];
  assign T196 = {T197, b3_real};
  assign T197 = T198 ? 21'h1fffff : 21'h0;
  assign T198 = b3_real[4'hf:4'hf];
  assign T199 = T200 ? 16'hffff : 16'h0;
  assign T200 = yz21_real[4'hf:4'hf];
  assign yz2_real = T205 + T201;
  assign T201 = T203 - T202;
  assign T202 = $signed(16'h1) * $signed(yz22_imag);
  assign T203 = $signed(16'h0) * $signed(T204);
  assign T204 = yz22_real + yz22_imag;
  assign T205 = {T206, yz21_real};
  assign T206 = T207 ? 16'hffff : 16'h0;
  assign T207 = yz21_real[4'hf:4'hf];
  assign yy3_imag = T208;
  assign T208 = T209[4'hf:1'h0];
  assign T209 = T27 ? yz3_imag : T210;
  assign T210 = T26 ? yz2_imag : yz3_imag;
  assign yz3_imag = T213 - T211;
  assign T211 = T168 + T212;
  assign T212 = $signed(16'h1) * $signed(yz22_real);
  assign T213 = {T231, yz21_imag};
  assign yz21_imag = T214;
  assign T214 = T215[4'hf:1'h0];
  assign T215 = T27 ? d2_imag : T216;
  assign T216 = T26 ? T228 : d2_imag;
  assign d2_imag = T217 + c5_imag;
  assign T217 = {T226, c2_imag};
  assign c2_imag = io_x0_imag - c22_imag;
  assign c22_imag = T218;
  assign T218 = T219[4'hf:1'h0];
  assign T219 = T193 ? T221 : T220;
  assign T220 = T192 ? T223 : T221;
  assign T221 = $signed(T222) / $signed(22'h100000);
  assign T222 = $signed(21'h80000) * $signed(b2_imag);
  assign T223 = {T224, io_x1_imag};
  assign T224 = T225 ? 21'h1fffff : 21'h0;
  assign T225 = io_x1_imag[4'hf:4'hf];
  assign T226 = T227 ? 21'h1fffff : 21'h0;
  assign T227 = c2_imag[4'hf:4'hf];
  assign T228 = {T229, b3_imag};
  assign T229 = T230 ? 21'h1fffff : 21'h0;
  assign T230 = b3_imag[4'hf:4'hf];
  assign T231 = T232 ? 16'hffff : 16'h0;
  assign T232 = yz21_imag[4'hf:4'hf];
  assign yz2_imag = T235 + T233;
  assign T233 = T203 + T234;
  assign T234 = $signed(16'h1) * $signed(yz22_real);
  assign T235 = {T236, yz21_imag};
  assign T236 = T237 ? 16'hffff : 16'h0;
  assign T237 = yz21_imag[4'hf:4'hf];
  assign T238 = $signed(yy3_real) * $signed(T239);
  assign T239 = io_twiddle3_real + io_twiddle3_imag;
  assign T240 = 4'h3 < io_radix;
  assign T241 = {T242, io_x3_imag};
  assign T242 = T243 ? 16'hffff : 16'h0;
  assign T243 = io_x3_imag[4'hf:4'hf];
  assign T244 = T240 == 1'h0;
  assign io_y3_real = T245;
  assign T245 = T246[4'hf:1'h0];
  assign T246 = T244 ? T253 : T247;
  assign T247 = T240 ? yx3_real : T248;
  assign T248 = {T249, io_x3_real};
  assign T249 = T250 ? 16'hffff : 16'h0;
  assign T250 = io_x3_real[4'hf:4'hf];
  assign yx3_real = T238 - T251;
  assign T251 = $signed(T252) * $signed(io_twiddle3_imag);
  assign T252 = yy3_real + yy3_imag;
  assign T253 = {T254, io_x3_real};
  assign T254 = T255 ? 16'hffff : 16'h0;
  assign T255 = io_x3_real[4'hf:4'hf];
  assign io_y2_imag = T256;
  assign T256 = T257[4'hf:1'h0];
  assign T257 = T296 ? T293 : T258;
  assign T258 = T292 ? yx2_imag : T259;
  assign T259 = {T260, io_x2_imag};
  assign T260 = T261 ? 16'hffff : 16'h0;
  assign T261 = io_x2_imag[4'hf:4'hf];
  assign yx2_imag = T290 + T262;
  assign T262 = $signed(T263) * $signed(io_twiddle2_real);
  assign T263 = yy2_imag - yy2_real;
  assign yy2_real = T264;
  assign T264 = T265[4'hf:1'h0];
  assign T265 = T22 ? T274 : T266;
  assign T266 = T19 ? T271 : T267;
  assign T267 = T18 ? yz4_real : T268;
  assign T268 = {T269, yz2_real};
  assign T269 = T270 ? 5'h1f : 5'h0;
  assign T270 = yz2_real[5'h1f:5'h1f];
  assign T271 = {T272, b5_real};
  assign T272 = T273 ? 21'h1fffff : 21'h0;
  assign T273 = b5_real[4'hf:4'hf];
  assign T274 = {T275, yz2_real};
  assign T275 = T276 ? 5'h1f : 5'h0;
  assign T276 = yz2_real[5'h1f:5'h1f];
  assign yy2_imag = T277;
  assign T277 = T278[4'hf:1'h0];
  assign T278 = T22 ? T287 : T279;
  assign T279 = T19 ? T284 : T280;
  assign T280 = T18 ? yz4_imag : T281;
  assign T281 = {T282, yz2_imag};
  assign T282 = T283 ? 5'h1f : 5'h0;
  assign T283 = yz2_imag[5'h1f:5'h1f];
  assign T284 = {T285, b5_imag};
  assign T285 = T286 ? 21'h1fffff : 21'h0;
  assign T286 = b5_imag[4'hf:4'hf];
  assign T287 = {T288, yz2_imag};
  assign T288 = T289 ? 5'h1f : 5'h0;
  assign T289 = yz2_imag[5'h1f:5'h1f];
  assign T290 = $signed(yy2_real) * $signed(T291);
  assign T291 = io_twiddle2_real + io_twiddle2_imag;
  assign T292 = 4'h2 < io_radix;
  assign T293 = {T294, io_x2_imag};
  assign T294 = T295 ? 16'hffff : 16'h0;
  assign T295 = io_x2_imag[4'hf:4'hf];
  assign T296 = T292 == 1'h0;
  assign io_y2_real = T297;
  assign T297 = T298[4'hf:1'h0];
  assign T298 = T296 ? T305 : T299;
  assign T299 = T292 ? yx2_real : T300;
  assign T300 = {T301, io_x2_real};
  assign T301 = T302 ? 16'hffff : 16'h0;
  assign T302 = io_x2_real[4'hf:4'hf];
  assign yx2_real = T290 - T303;
  assign T303 = $signed(T304) * $signed(io_twiddle2_imag);
  assign T304 = yy2_real + yy2_imag;
  assign T305 = {T306, io_x2_real};
  assign T306 = T307 ? 16'hffff : 16'h0;
  assign T307 = io_x2_real[4'hf:4'hf];
  assign io_y1_imag = T308;
  assign T308 = T309[4'hf:1'h0];
  assign T309 = T346 + T310;
  assign T310 = $signed(T311) * $signed(io_twiddle1_real);
  assign T311 = yy1_imag - yy1_real;
  assign yy1_real = T312;
  assign T312 = T313[4'hf:1'h0];
  assign T313 = T90 ? yz1_real : T314;
  assign T314 = T86 ? T327 : T315;
  assign T315 = T83 ? yz1_real : T316;
  assign T316 = T82 ? T324 : yz1_real;
  assign yz1_real = d1_real + T317;
  assign T317 = {T322, T318};
  assign T318 = T320 - T319;
  assign T319 = $signed(16'h1) * $signed(d4_imag);
  assign T320 = $signed(16'h0) * $signed(T321);
  assign T321 = d4_real + d4_imag;
  assign T322 = T323 ? 5'h1f : 5'h0;
  assign T323 = T318[5'h1f:5'h1f];
  assign T324 = {T325, c2_real};
  assign T325 = T326 ? 21'h1fffff : 21'h0;
  assign T326 = c2_real[4'hf:4'hf];
  assign T327 = {T328, yz3_real};
  assign T328 = T329 ? 5'h1f : 5'h0;
  assign T329 = yz3_real[5'h1f:5'h1f];
  assign yy1_imag = T330;
  assign T330 = T331[4'hf:1'h0];
  assign T331 = T90 ? yz1_imag : T332;
  assign T332 = T86 ? T343 : T333;
  assign T333 = T83 ? yz1_imag : T334;
  assign T334 = T82 ? T340 : yz1_imag;
  assign yz1_imag = d1_imag + T335;
  assign T335 = {T338, T336};
  assign T336 = T320 + T337;
  assign T337 = $signed(16'h1) * $signed(d4_real);
  assign T338 = T339 ? 5'h1f : 5'h0;
  assign T339 = T336[5'h1f:5'h1f];
  assign T340 = {T341, c2_imag};
  assign T341 = T342 ? 21'h1fffff : 21'h0;
  assign T342 = c2_imag[4'hf:4'hf];
  assign T343 = {T344, yz3_imag};
  assign T344 = T345 ? 5'h1f : 5'h0;
  assign T345 = yz3_imag[5'h1f:5'h1f];
  assign T346 = $signed(yy1_real) * $signed(T347);
  assign T347 = io_twiddle1_real + io_twiddle1_imag;
  assign io_y1_real = T348;
  assign T348 = T349[4'hf:1'h0];
  assign T349 = T346 - T350;
  assign T350 = $signed(T351) * $signed(io_twiddle1_imag);
  assign T351 = yy1_real + yy1_imag;
  assign io_y0_imag = T352;
  assign T352 = T90 ? yz0_imag : T353;
  assign T353 = T86 ? c7_imag : T354;
  assign T354 = T83 ? yz0_imag : T355;
  assign T355 = T82 ? b1_imag : yz0_imag;
  assign yz0_imag = io_x0_imag + d02_imag;
  assign d02_imag = T356;
  assign T356 = T31 ? c7_imag : T357;
  assign T357 = T30 ? b1_imag : c7_imag;
  assign c7_imag = b1_imag + b2_imag;
  assign io_y0_real = T358;
  assign T358 = T90 ? yz0_real : T359;
  assign T359 = T86 ? c7_real : T360;
  assign T360 = T83 ? yz0_real : T361;
  assign T361 = T82 ? b1_real : yz0_real;
  assign yz0_real = io_x0_real + d02_real;
  assign d02_real = T362;
  assign T362 = T31 ? c7_real : T363;
  assign T363 = T30 ? b1_real : c7_real;
  assign c7_real = b1_real + b2_real;
endmodule

